module fc2 (
	input [127:0] in,
	output [127:0] out
);

wire [3:0] relu_out [0:31];
wire [8:0] weighted_sum [0:31];
wire [8:0] sharing0;
wire [8:0] sharing1;
wire [8:0] sharing2;
wire [8:0] sharing3;
wire [8:0] sharing4;
wire [8:0] sharing5;
wire [8:0] sharing6;
wire [8:0] sharing7;
wire [8:0] sharing8;
wire [8:0] sharing9;
wire [8:0] sharing10;
wire [8:0] sharing11;
wire [8:0] sharing12;
wire [8:0] sharing13;
wire [8:0] sharing14;
wire [8:0] sharing15;
wire [8:0] sharing16;
wire [8:0] sharing17;
wire [8:0] sharing18;
wire [8:0] sharing19;
wire [8:0] sharing20;
wire [8:0] sharing21;
wire [8:0] sharing22;
wire [8:0] sharing23;
wire [8:0] sharing24;
wire [8:0] sharing25;
wire [8:0] sharing26;
wire [8:0] sharing27;
wire [8:0] sharing28;
wire [8:0] sharing29;
wire [8:0] sharing30;
wire [8:0] sharing31;
wire [8:0] sharing32;
wire [8:0] sharing33;
wire [8:0] sharing34;
wire [8:0] sharing35;
wire [8:0] sharing36;
wire [8:0] sharing37;
wire [8:0] sharing38;
wire [8:0] sharing39;
wire [8:0] sharing40;
wire [8:0] sharing41;
wire [8:0] sharing42;
wire [8:0] sharing43;
wire [8:0] sharing44;
wire [8:0] sharing45;
wire [8:0] sharing46;
wire [8:0] sharing47;
wire [8:0] sharing48;
wire [8:0] sharing49;

assign sharing0 = $signed(in[123-:4])+$signed(-in[107-:4])+$signed(-in[103-:4]);
assign sharing1 = $signed({in[71-:4],1'b0})+$signed({in[31-:4],1'b0})+$signed(-{in[91-:4],1'b0})+$signed(-in[43-:4])+$signed(-in[7-:4])+$signed(-in[127-:4]);
assign sharing2 = $signed(in[103-:4])+$signed(in[11-:4])+$signed({in[15-:4],1'b0})+$signed(in[79-:4])+$signed({in[19-:4],1'b0})+$signed(in[87-:4])+$signed(-{in[87-:4],2'b0})+$signed(-{in[71-:4],1'b0});
assign sharing3 = $signed(in[67-:4])+$signed({in[43-:4],1'b0})+$signed(in[75-:4])+$signed(in[119-:4])+$signed(-{in[107-:4],1'b0})+$signed(-in[47-:4])+$signed(-in[115-:4])+$signed(-in[23-:4])+$signed(-{in[27-:4],2'b0});
assign sharing4 = $signed(in[3-:4])+$signed(in[55-:4])+$signed(-in[35-:4])+$signed(-in[27-:4])+$signed(-in[23-:4])+$signed(-in[119-:4]);
assign sharing5 = $signed({in[75-:4],1'b0})+$signed(in[43-:4])+$signed({in[59-:4],1'b0})+$signed(in[15-:4])+$signed(-{in[95-:4],1'b0})+$signed(-in[47-:4]);
assign sharing6 = $signed(in[75-:4])+$signed(in[107-:4])+$signed(in[15-:4])+$signed(in[95-:4])+$signed(in[31-:4])+$signed(-{in[39-:4],1'b0})+$signed(-{in[107-:4],2'b0})+$signed(-in[115-:4])+$signed(-in[35-:4]);
assign sharing7 = $signed(in[43-:4])+$signed(in[11-:4])+$signed({in[87-:4],1'b0})+$signed(-in[99-:4])+$signed(-{in[71-:4],1'b0})+$signed(-in[103-:4])+$signed(-{in[47-:4],1'b0})+$signed(-{in[59-:4],1'b0})+$signed(-in[27-:4])+$signed(-in[127-:4]);
assign sharing8 = $signed({in[99-:4],1'b0})+$signed({in[43-:4],1'b0})+$signed(in[11-:4])+$signed(in[47-:4])+$signed(in[55-:4])+$signed({in[95-:4],1'b0})+$signed(-in[35-:4])+$signed(-{in[83-:4],1'b0})+$signed(-in[91-:4]);
assign sharing9 = $signed({in[103-:4],1'b0})+$signed(in[39-:4])+$signed(in[7-:4])+$signed(in[15-:4])+$signed(in[115-:4])+$signed(in[31-:4])+$signed(-in[123-:4])+$signed(-in[71-:4]);
assign sharing10 = $signed(in[123-:4])+$signed({in[123-:4],1'b0})+$signed(in[91-:4])+$signed(in[71-:4])+$signed(-in[19-:4])+$signed(-in[63-:4]);
assign sharing11 = $signed({in[79-:4],1'b0})+$signed(in[15-:4])+$signed(-in[7-:4])+$signed(-in[103-:4])+$signed(-{in[75-:4],1'b0})+$signed(-{in[47-:4],1'b0})+$signed(-{in[27-:4],1'b0});
assign sharing12 = $signed(-{in[103-:4],1'b0})+$signed(-in[59-:4])+$signed(-in[107-:4])+$signed(-in[75-:4])+$signed(-in[47-:4])+$signed(-in[15-:4])+$signed(-in[51-:4])+$signed(-in[119-:4])+$signed(-in[23-:4])+$signed(-in[27-:4])+$signed(-in[127-:4]);
assign sharing13 = $signed(in[3-:4])+$signed(in[39-:4])+$signed(in[75-:4])+$signed(in[79-:4])+$signed({in[51-:4],1'b0})+$signed(in[51-:4])+$signed({in[115-:4],1'b0})+$signed({in[27-:4],1'b0})+$signed({in[63-:4],1'b0})+$signed(-in[43-:4])+$signed(-in[83-:4])+$signed(-{in[47-:4],1'b0});
assign sharing14 = $signed(in[59-:4])+$signed(-in[91-:4])+$signed(-in[19-:4])+$signed(-in[127-:4]);
assign sharing15 = $signed(in[115-:4])+$signed(in[51-:4])+$signed({in[55-:4],1'b0})+$signed(in[71-:4])+$signed(-{in[123-:4],1'b0});
assign sharing16 = $signed({in[3-:4],1'b0})+$signed(-{in[99-:4],1'b0})+$signed(-in[39-:4])+$signed(-in[79-:4])+$signed(-{in[127-:4],1'b0})+$signed(-in[63-:4]);
assign sharing17 = $signed({in[3-:4],1'b0})+$signed(in[55-:4])+$signed(in[95-:4])+$signed(in[63-:4])+$signed(-in[67-:4])+$signed(-in[99-:4]);
assign sharing18 = $signed(in[27-:4])+$signed({in[111-:4],1'b0})+$signed(in[31-:4])+$signed(-{in[83-:4],1'b0})+$signed(-{in[103-:4],1'b0})+$signed(-{in[115-:4],1'b0});
assign sharing19 = $signed({in[67-:4],1'b0})+$signed({in[103-:4],1'b0})+$signed(in[11-:4])+$signed({in[83-:4],1'b0})+$signed(in[23-:4])+$signed(in[31-:4])+$signed(-{in[115-:4],1'b0})+$signed(-in[123-:4]);
assign sharing20 = $signed({in[119-:4],1'b0})+$signed(in[55-:4])+$signed(-{in[75-:4],1'b0})+$signed(-in[71-:4])+$signed(-{in[111-:4],1'b0})+$signed(-in[95-:4]);
assign sharing21 = $signed({in[39-:4],1'b0})+$signed(in[71-:4])+$signed(in[103-:4])+$signed(in[15-:4])+$signed({in[83-:4],1'b0})+$signed(in[83-:4])+$signed(-in[35-:4])+$signed(-{in[51-:4],1'b0})+$signed(-in[19-:4])+$signed(-in[127-:4])+$signed(-in[63-:4]);
assign sharing22 = $signed(in[7-:4])+$signed(in[75-:4])+$signed(in[79-:4])+$signed(in[119-:4])+$signed(in[27-:4])+$signed(-in[11-:4]);
assign sharing23 = $signed({in[11-:4],1'b0})+$signed(in[11-:4])+$signed(in[111-:4])+$signed({in[51-:4],1'b0})+$signed(in[91-:4])+$signed(in[127-:4])+$signed(-{in[71-:4],1'b0});
assign sharing24 = $signed({in[15-:4],1'b0})+$signed(in[31-:4])+$signed(-in[3-:4])+$signed(-in[87-:4]);
assign sharing25 = $signed({in[35-:4],1'b0})+$signed(in[67-:4])+$signed(in[99-:4])+$signed(in[107-:4])+$signed(in[111-:4])+$signed({in[115-:4],1'b0})+$signed({in[119-:4],1'b0})+$signed(-{in[11-:4],1'b0})+$signed(-in[59-:4])+$signed(-{in[43-:4],1'b0})+$signed(-{in[127-:4],2'b0});
assign sharing26 = $signed({in[3-:4],1'b0})+$signed(in[123-:4])+$signed(-in[91-:4])+$signed(-in[7-:4]);
assign sharing27 = $signed(in[3-:4])+$signed(in[35-:4])+$signed(in[75-:4])+$signed({in[111-:4],1'b0})+$signed({in[19-:4],2'b0})+$signed(in[51-:4])+$signed({in[95-:4],1'b0})+$signed(in[63-:4])+$signed(-{in[39-:4],1'b0})+$signed(-in[27-:4])+$signed(-{in[103-:4],1'b0})+$signed(-in[55-:4]);
assign sharing28 = $signed({in[23-:4],1'b0})+$signed(-in[43-:4])+$signed(-in[115-:4])+$signed(-in[87-:4])+$signed(-in[127-:4]);
assign sharing29 = $signed({in[43-:4],1'b0})+$signed(in[75-:4])+$signed(in[79-:4])+$signed(in[47-:4])+$signed(in[19-:4])+$signed({in[91-:4],1'b0})+$signed(-in[127-:4])+$signed(-in[95-:4]);
assign sharing30 = $signed(in[3-:4])+$signed(in[99-:4])+$signed(-in[39-:4])+$signed(-{in[51-:4],1'b0})+$signed(-in[115-:4])+$signed(-in[87-:4])+$signed(-in[123-:4])+$signed(-{in[63-:4],1'b0});
assign sharing31 = $signed(in[75-:4])+$signed({in[87-:4],1'b0})+$signed({in[15-:4],1'b0});
assign sharing32 = $signed(in[99-:4])+$signed(-in[83-:4])+$signed(-{in[115-:4],1'b0})+$signed(-in[123-:4])+$signed(-in[7-:4]);
assign sharing33 = $signed({in[23-:4],1'b0})+$signed(in[111-:4])+$signed(-{in[27-:4],3'b0})+$signed(-in[91-:4]);
assign sharing34 = $signed({in[127-:4],1'b0})+$signed(in[39-:4])+$signed(-{in[59-:4],1'b0})+$signed(-{in[87-:4],2'b0});
assign sharing35 = $signed({in[111-:4],1'b0})+$signed({in[59-:4],1'b0})+$signed(in[27-:4])+$signed(in[63-:4])+$signed(in[95-:4])+$signed(-{in[63-:4],2'b0});
assign sharing36 = $signed(in[107-:4])+$signed(in[59-:4])+$signed(-in[3-:4]);
assign sharing37 = $signed(in[47-:4])+$signed(-{in[87-:4],1'b0})+$signed(-in[111-:4]);
assign sharing38 = $signed(in[59-:4])+$signed(in[51-:4])+$signed({in[39-:4],1'b0})+$signed(-{in[47-:4],2'b0});
assign sharing39 = $signed({in[35-:4],1'b0})+$signed(in[83-:4])+$signed(-{in[107-:4],1'b0});
assign sharing40 = $signed(in[51-:4])+$signed(in[111-:4])+$signed(-in[83-:4])+$signed(-in[7-:4]);
assign sharing41 = $signed(in[63-:4])+$signed(-in[79-:4])+$signed(-{in[71-:4],1'b0})+$signed(-in[31-:4]);
assign sharing42 = $signed({in[35-:4],2'b0})+$signed({in[11-:4],1'b0})+$signed(in[115-:4]);
assign sharing43 = $signed({in[99-:4],2'b0})+$signed(-in[59-:4])+$signed(-{in[87-:4],1'b0});
assign sharing44 = $signed({in[71-:4],1'b0})+$signed({in[31-:4],1'b0})+$signed(-{in[111-:4],1'b0})+$signed(-in[23-:4]);
assign sharing45 = $signed({in[67-:4],1'b0})+$signed(in[75-:4])+$signed(-{in[95-:4],1'b0});
assign sharing46 = $signed({in[19-:4],1'b0})+$signed(in[87-:4])+$signed(-{in[39-:4],1'b0});
assign sharing47 = $signed({in[23-:4],2'b0})+$signed({in[87-:4],1'b0})+$signed(-{in[127-:4],2'b0});
assign sharing48 = $signed({in[27-:4],1'b0})+$signed(in[99-:4])+$signed(-{in[23-:4],1'b0});
assign sharing49 = $signed({in[59-:4],1'b0})+$signed({in[107-:4],1'b0})+$signed(in[31-:4]);
assign weighted_sum[0] = $signed(-in[99-:4])+$signed(-{in[27-:4],1'b0})+$signed(in[75-:4])+$signed({in[15-:4],1'b0})+$signed(-in[79-:4])+$signed({in[19-:4],2'b0})+$signed(-in[87-:4])+$signed(-{in[59-:4],1'b0})+$signed(-{in[63-:4],3'b0})+$signed({in[63-:4],1'b0})+$signed(sharing0)+$signed(sharing1)+$signed(sharing42)+$signed(1);
assign weighted_sum[1] = $signed(in[35-:4])+$signed({in[7-:4],1'b0})+$signed(-{in[43-:4],2'b0})+$signed(-{in[79-:4],1'b0})+$signed(-{in[51-:4],1'b0})+$signed(in[115-:4])+$signed({in[55-:4],1'b0})+$signed({in[91-:4],1'b0})+$signed(-{in[63-:4],2'b0})+$signed(-in[127-:4])+$signed(sharing17)+$signed(-sharing18)+$signed(sharing31)+$signed(-2);
assign weighted_sum[2] = $signed(-{in[35-:4],2'b0})+$signed(in[35-:4])+$signed(-{in[11-:4],2'b0})+$signed(in[59-:4])+$signed(-{in[51-:4],2'b0})+$signed(-{in[59-:4],3'b0})+$signed({in[91-:4],1'b0})+$signed(-in[123-:4])+$signed(-{in[31-:4],2'b0})+$signed(sharing2)+$signed(sharing3)+$signed(sharing35)+$signed(-4);
assign weighted_sum[3] = $signed({in[3-:4],2'b0})+$signed(-in[67-:4])+$signed({in[103-:4],2'b0})+$signed({in[7-:4],1'b0})+$signed(-in[111-:4])+$signed({in[83-:4],2'b0})+$signed(-in[19-:4])+$signed(-{in[55-:4],2'b0})+$signed(-{in[123-:4],1'b0})+$signed(in[59-:4])+$signed({in[127-:4],2'b0})+$signed({in[63-:4],1'b0})+$signed(sharing4)+$signed(sharing5)+$signed(0);
assign weighted_sum[4] = $signed({in[3-:4],1'b0})+$signed({in[7-:4],2'b0})+$signed(in[91-:4])+$signed({in[111-:4],1'b0})+$signed(in[79-:4])+$signed(-{in[55-:4],1'b0})+$signed(in[119-:4])+$signed(-in[123-:4])+$signed(in[63-:4])+$signed(sharing6)+$signed(sharing7)+$signed(-4);
assign weighted_sum[5] = $signed({in[39-:4],1'b0})+$signed(-{in[75-:4],2'b0})+$signed(-{in[111-:4],3'b0})+$signed({in[79-:4],1'b0})+$signed(in[27-:4])+$signed(-in[63-:4])+$signed(-in[95-:4])+$signed(in[127-:4])+$signed(sharing25)+$signed(-sharing26)+$signed(sharing31)+$signed(-sharing44)+$signed(2);
assign weighted_sum[6] = $signed({in[11-:4],1'b0})+$signed(-{in[107-:4],1'b0})+$signed(in[115-:4])+$signed(-in[51-:4])+$signed({in[55-:4],1'b0})+$signed({in[91-:4],2'b0})+$signed(in[127-:4])+$signed(sharing4)+$signed(-sharing5)+$signed(-sharing32)+$signed(sharing41)+$signed(-sharing46)+$signed(-3);
assign weighted_sum[7] = $signed({in[35-:4],1'b0})+$signed({in[99-:4],1'b0})+$signed(in[103-:4])+$signed(-in[27-:4])+$signed({in[51-:4],1'b0})+$signed(-in[19-:4])+$signed({in[31-:4],1'b0})+$signed(-{in[91-:4],2'b0})+$signed(in[91-:4])+$signed(-{in[95-:4],2'b0})+$signed({in[63-:4],1'b0})+$signed(sharing19)+$signed(-sharing20)+$signed(sharing36)+$signed(-sharing37)+$signed(1);
assign weighted_sum[8] = $signed(-{in[3-:4],2'b0})+$signed({in[11-:4],1'b0})+$signed(in[75-:4])+$signed({in[111-:4],2'b0})+$signed(-{in[15-:4],2'b0})+$signed({in[51-:4],1'b0})+$signed(-in[19-:4])+$signed({in[115-:4],1'b0})+$signed(in[23-:4])+$signed(-{in[31-:4],2'b0})+$signed({in[127-:4],1'b0})+$signed(sharing8)+$signed(sharing9)+$signed(sharing43)+$signed(2);
assign weighted_sum[9] = $signed({in[99-:4],1'b0})+$signed(in[99-:4])+$signed(in[107-:4])+$signed(in[111-:4])+$signed(-{in[115-:4],1'b0})+$signed({in[23-:4],2'b0})+$signed(-in[87-:4])+$signed(in[119-:4])+$signed({in[59-:4],2'b0})+$signed({in[91-:4],1'b0})+$signed({in[31-:4],2'b0})+$signed(in[95-:4])+$signed(sharing10)+$signed(sharing11)+$signed(-2);
assign weighted_sum[10] = $signed(in[67-:4])+$signed(in[43-:4])+$signed(-in[111-:4])+$signed(-in[87-:4])+$signed(-in[91-:4])+$signed(sharing12)+$signed(sharing32)+$signed(-2);
assign weighted_sum[11] = $signed({in[123-:4],1'b0})+$signed(-in[43-:4])+$signed(in[55-:4])+$signed(-in[87-:4])+$signed(sharing21)+$signed(-sharing22)+$signed(sharing44)+$signed(sharing49)+$signed(-2);
assign weighted_sum[12] = $signed(-{in[99-:4],1'b0})+$signed(in[35-:4])+$signed(in[27-:4])+$signed(-{in[79-:4],2'b0})+$signed(in[15-:4])+$signed(-{in[23-:4],1'b0})+$signed(-in[55-:4])+$signed(-in[123-:4])+$signed(in[95-:4])+$signed(sharing13)+$signed(sharing14)+$signed(sharing42)+$signed(sharing49)+$signed(3);
assign weighted_sum[13] = $signed(in[35-:4])+$signed(-{in[11-:4],2'b0})+$signed(in[107-:4])+$signed(-in[43-:4])+$signed({in[111-:4],1'b0})+$signed(-in[47-:4])+$signed(-{in[51-:4],2'b0})+$signed({in[115-:4],1'b0})+$signed(in[83-:4])+$signed(in[119-:4])+$signed({in[27-:4],1'b0})+$signed(sharing15)+$signed(sharing16)+$signed(sharing33)+$signed(sharing45)+$signed(-2);
assign weighted_sum[14] = $signed(-{in[71-:4],2'b0})+$signed({in[103-:4],1'b0})+$signed(in[71-:4])+$signed(-{in[75-:4],2'b0})+$signed(-{in[15-:4],2'b0})+$signed({in[111-:4],1'b0})+$signed(in[15-:4])+$signed(-{in[19-:4],2'b0})+$signed({in[23-:4],1'b0})+$signed(-in[119-:4])+$signed({in[87-:4],1'b0})+$signed({in[27-:4],1'b0})+$signed(-in[59-:4])+$signed(-in[31-:4])+$signed(sharing29)+$signed(-sharing30)+$signed(0);
assign weighted_sum[15] = $signed(in[3-:4])+$signed({in[7-:4],1'b0})+$signed(-{in[47-:4],3'b0})+$signed({in[83-:4],1'b0})+$signed(-in[19-:4])+$signed(in[23-:4])+$signed(-{in[23-:4],2'b0})+$signed(-in[55-:4])+$signed({in[91-:4],1'b0})+$signed(sharing6)+$signed(-sharing7)+$signed(-sharing40)+$signed(0);
assign weighted_sum[16] = $signed(in[3-:4])+$signed(-{in[7-:4],2'b0})+$signed(in[7-:4])+$signed(-in[107-:4])+$signed(in[47-:4])+$signed(in[79-:4])+$signed(-in[51-:4])+$signed(sharing17)+$signed(sharing18)+$signed(sharing33)+$signed(sharing46)+$signed(0);
assign weighted_sum[17] = $signed(-{in[3-:4],2'b0})+$signed({in[103-:4],1'b0})+$signed({in[7-:4],1'b0})+$signed({in[43-:4],1'b0})+$signed(-in[107-:4])+$signed(in[115-:4])+$signed(-{in[119-:4],1'b0})+$signed(-in[23-:4])+$signed(in[63-:4])+$signed(sharing23)+$signed(-sharing24)+$signed(sharing34)+$signed(-1);
assign weighted_sum[18] = $signed(-{in[67-:4],2'b0})+$signed(in[3-:4])+$signed(-in[79-:4])+$signed({in[19-:4],1'b0})+$signed({in[123-:4],1'b0})+$signed({in[127-:4],2'b0})+$signed(sharing8)+$signed(-sharing9)+$signed(sharing35)+$signed(2);
assign weighted_sum[19] = $signed(-in[11-:4])+$signed(-in[43-:4])+$signed(-in[19-:4])+$signed(-{in[55-:4],1'b0})+$signed(-{in[91-:4],1'b0})+$signed(sharing12)+$signed(sharing41)+$signed(-2);
assign weighted_sum[20] = $signed({in[67-:4],2'b0})+$signed({in[35-:4],1'b0})+$signed(in[99-:4])+$signed(-{in[99-:4],2'b0})+$signed(-{in[71-:4],2'b0})+$signed(in[71-:4])+$signed(-in[11-:4])+$signed({in[15-:4],2'b0})+$signed(in[111-:4])+$signed({in[119-:4],1'b0})+$signed({in[91-:4],1'b0})+$signed(-{in[31-:4],1'b0})+$signed(sharing13)+$signed(-sharing14)+$signed(sharing47)+$signed(-2);
assign weighted_sum[21] = $signed({in[91-:4],2'b0})+$signed(-{in[35-:4],1'b0})+$signed({in[43-:4],1'b0})+$signed(-{in[75-:4],1'b0})+$signed({in[111-:4],1'b0})+$signed(in[47-:4])+$signed({in[19-:4],1'b0})+$signed({in[119-:4],2'b0})+$signed(-{in[123-:4],2'b0})+$signed(in[27-:4])+$signed({in[95-:4],1'b0})+$signed(sharing0)+$signed(-sharing1)+$signed(sharing38)+$signed(sharing47)+$signed(-1);
assign weighted_sum[22] = $signed(-{in[7-:4],1'b0})+$signed({in[39-:4],1'b0})+$signed(in[39-:4])+$signed({in[107-:4],2'b0})+$signed(in[43-:4])+$signed({in[79-:4],2'b0})+$signed({in[15-:4],1'b0})+$signed(-{in[51-:4],2'b0})+$signed(in[51-:4])+$signed(-{in[55-:4],2'b0})+$signed(in[119-:4])+$signed({in[59-:4],1'b0})+$signed(-in[127-:4])+$signed(sharing19)+$signed(sharing20)+$signed(-sharing48)+$signed(2);
assign weighted_sum[23] = $signed(-{in[35-:4],1'b0})+$signed(-in[3-:4])+$signed(in[43-:4])+$signed({in[51-:4],1'b0})+$signed(-{in[119-:4],1'b0})+$signed(-in[23-:4])+$signed(-{in[123-:4],3'b0})+$signed(in[27-:4])+$signed(in[31-:4])+$signed(sharing10)+$signed(-sharing11)+$signed(-sharing34)+$signed(sharing45)+$signed(0);
assign weighted_sum[24] = $signed(in[67-:4])+$signed(-{in[71-:4],2'b0})+$signed({in[103-:4],1'b0})+$signed(-{in[43-:4],1'b0})+$signed({in[15-:4],1'b0})+$signed({in[119-:4],1'b0})+$signed(-{in[27-:4],2'b0})+$signed(in[123-:4])+$signed(-{in[59-:4],2'b0})+$signed(-in[95-:4])+$signed(sharing21)+$signed(sharing22)+$signed(sharing36)+$signed(sharing37)+$signed(0);
assign weighted_sum[25] = $signed({in[35-:4],1'b0})+$signed(in[103-:4])+$signed(-{in[107-:4],1'b0})+$signed(in[43-:4])+$signed(-in[75-:4])+$signed({in[83-:4],1'b0})+$signed(-{in[119-:4],2'b0})+$signed(-{in[55-:4],1'b0})+$signed(in[123-:4])+$signed({in[63-:4],2'b0})+$signed(sharing23)+$signed(sharing24)+$signed(sharing38)+$signed(sharing48)+$signed(0);
assign weighted_sum[26] = $signed(-{in[99-:4],2'b0})+$signed({in[67-:4],1'b0})+$signed(in[103-:4])+$signed(-in[71-:4])+$signed(in[39-:4])+$signed({in[15-:4],2'b0})+$signed(-in[79-:4])+$signed(in[19-:4])+$signed(in[115-:4])+$signed(-{in[23-:4],1'b0})+$signed(in[55-:4])+$signed(-in[87-:4])+$signed(sharing25)+$signed(sharing26)+$signed(1);
assign weighted_sum[27] = $signed(in[91-:4])+$signed(in[11-:4])+$signed(-{in[79-:4],1'b0})+$signed({in[15-:4],1'b0})+$signed(-in[47-:4])+$signed(-{in[83-:4],2'b0})+$signed(in[19-:4])+$signed({in[119-:4],1'b0})+$signed({in[59-:4],1'b0})+$signed(-in[123-:4])+$signed(in[31-:4])+$signed(-{in[63-:4],2'b0})+$signed({in[31-:4],1'b0})+$signed(in[95-:4])+$signed(sharing27)+$signed(sharing28)+$signed(sharing39)+$signed(2);
assign weighted_sum[28] = $signed({in[35-:4],1'b0})+$signed(-{in[103-:4],2'b0})+$signed(-{in[111-:4],2'b0})+$signed({in[79-:4],1'b0})+$signed({in[51-:4],1'b0})+$signed(-in[55-:4])+$signed(-{in[63-:4],1'b0})+$signed({in[95-:4],1'b0})+$signed({in[123-:4],1'b0})+$signed(-{in[127-:4],1'b0})+$signed(sharing2)+$signed(-sharing3)+$signed(sharing40)+$signed(2);
assign weighted_sum[29] = $signed(in[67-:4])+$signed(in[103-:4])+$signed(-in[7-:4])+$signed(-{in[11-:4],2'b0})+$signed({in[75-:4],1'b0})+$signed(in[11-:4])+$signed({in[111-:4],2'b0})+$signed({in[119-:4],2'b0})+$signed(-{in[91-:4],3'b0})+$signed(in[91-:4])+$signed(sharing29)+$signed(sharing30)+$signed(-sharing39)+$signed(3);
assign weighted_sum[30] = $signed({in[35-:4],2'b0})+$signed(-{in[67-:4],1'b0})+$signed({in[91-:4],1'b0})+$signed(-{in[71-:4],1'b0})+$signed(-in[107-:4])+$signed({in[47-:4],1'b0})+$signed(in[119-:4])+$signed(-{in[59-:4],2'b0})+$signed({in[123-:4],1'b0})+$signed({in[127-:4],1'b0})+$signed(sharing27)+$signed(-sharing28)+$signed(-sharing43)+$signed(0);
assign weighted_sum[31] = $signed(-{in[67-:4],2'b0})+$signed(in[67-:4])+$signed({in[7-:4],1'b0})+$signed(in[103-:4])+$signed({in[75-:4],1'b0})+$signed({in[107-:4],1'b0})+$signed(-{in[79-:4],2'b0})+$signed({in[47-:4],1'b0})+$signed({in[115-:4],2'b0})+$signed(in[19-:4])+$signed(-{in[63-:4],3'b0})+$signed({in[63-:4],1'b0})+$signed(in[95-:4])+$signed(sharing15)+$signed(-sharing16)+$signed(1);
assign relu_out[0] = (weighted_sum[0][8]==1) ? 4'd0 : (weighted_sum[0][7:3] > 6 ? 4'd6 : weighted_sum[0][6:3]);
assign relu_out[1] = (weighted_sum[1][8]==1) ? 4'd0 : (weighted_sum[1][7:3] > 6 ? 4'd6 : weighted_sum[1][6:3]);
assign relu_out[2] = (weighted_sum[2][8]==1) ? 4'd0 : (weighted_sum[2][7:3] > 6 ? 4'd6 : weighted_sum[2][6:3]);
assign relu_out[3] = (weighted_sum[3][8]==1) ? 4'd0 : (weighted_sum[3][7:3] > 6 ? 4'd6 : weighted_sum[3][6:3]);
assign relu_out[4] = (weighted_sum[4][8]==1) ? 4'd0 : (weighted_sum[4][7:3] > 6 ? 4'd6 : weighted_sum[4][6:3]);
assign relu_out[5] = (weighted_sum[5][8]==1) ? 4'd0 : (weighted_sum[5][7:3] > 6 ? 4'd6 : weighted_sum[5][6:3]);
assign relu_out[6] = (weighted_sum[6][8]==1) ? 4'd0 : (weighted_sum[6][7:3] > 6 ? 4'd6 : weighted_sum[6][6:3]);
assign relu_out[7] = (weighted_sum[7][8]==1) ? 4'd0 : (weighted_sum[7][7:3] > 6 ? 4'd6 : weighted_sum[7][6:3]);
assign relu_out[8] = (weighted_sum[8][8]==1) ? 4'd0 : (weighted_sum[8][7:3] > 6 ? 4'd6 : weighted_sum[8][6:3]);
assign relu_out[9] = (weighted_sum[9][8]==1) ? 4'd0 : (weighted_sum[9][7:3] > 6 ? 4'd6 : weighted_sum[9][6:3]);
assign relu_out[10] = (weighted_sum[10][8]==1) ? 4'd0 : (weighted_sum[10][7:3] > 6 ? 4'd6 : weighted_sum[10][6:3]);
assign relu_out[11] = (weighted_sum[11][8]==1) ? 4'd0 : (weighted_sum[11][7:3] > 6 ? 4'd6 : weighted_sum[11][6:3]);
assign relu_out[12] = (weighted_sum[12][8]==1) ? 4'd0 : (weighted_sum[12][7:3] > 6 ? 4'd6 : weighted_sum[12][6:3]);
assign relu_out[13] = (weighted_sum[13][8]==1) ? 4'd0 : (weighted_sum[13][7:3] > 6 ? 4'd6 : weighted_sum[13][6:3]);
assign relu_out[14] = (weighted_sum[14][8]==1) ? 4'd0 : (weighted_sum[14][7:3] > 6 ? 4'd6 : weighted_sum[14][6:3]);
assign relu_out[15] = (weighted_sum[15][8]==1) ? 4'd0 : (weighted_sum[15][7:3] > 6 ? 4'd6 : weighted_sum[15][6:3]);
assign relu_out[16] = (weighted_sum[16][8]==1) ? 4'd0 : (weighted_sum[16][7:3] > 6 ? 4'd6 : weighted_sum[16][6:3]);
assign relu_out[17] = (weighted_sum[17][8]==1) ? 4'd0 : (weighted_sum[17][7:3] > 6 ? 4'd6 : weighted_sum[17][6:3]);
assign relu_out[18] = (weighted_sum[18][8]==1) ? 4'd0 : (weighted_sum[18][7:3] > 6 ? 4'd6 : weighted_sum[18][6:3]);
assign relu_out[19] = (weighted_sum[19][8]==1) ? 4'd0 : (weighted_sum[19][7:3] > 6 ? 4'd6 : weighted_sum[19][6:3]);
assign relu_out[20] = (weighted_sum[20][8]==1) ? 4'd0 : (weighted_sum[20][7:3] > 6 ? 4'd6 : weighted_sum[20][6:3]);
assign relu_out[21] = (weighted_sum[21][8]==1) ? 4'd0 : (weighted_sum[21][7:3] > 6 ? 4'd6 : weighted_sum[21][6:3]);
assign relu_out[22] = (weighted_sum[22][8]==1) ? 4'd0 : (weighted_sum[22][7:3] > 6 ? 4'd6 : weighted_sum[22][6:3]);
assign relu_out[23] = (weighted_sum[23][8]==1) ? 4'd0 : (weighted_sum[23][7:3] > 6 ? 4'd6 : weighted_sum[23][6:3]);
assign relu_out[24] = (weighted_sum[24][8]==1) ? 4'd0 : (weighted_sum[24][7:3] > 6 ? 4'd6 : weighted_sum[24][6:3]);
assign relu_out[25] = (weighted_sum[25][8]==1) ? 4'd0 : (weighted_sum[25][7:3] > 6 ? 4'd6 : weighted_sum[25][6:3]);
assign relu_out[26] = (weighted_sum[26][8]==1) ? 4'd0 : (weighted_sum[26][7:3] > 6 ? 4'd6 : weighted_sum[26][6:3]);
assign relu_out[27] = (weighted_sum[27][8]==1) ? 4'd0 : (weighted_sum[27][7:3] > 6 ? 4'd6 : weighted_sum[27][6:3]);
assign relu_out[28] = (weighted_sum[28][8]==1) ? 4'd0 : (weighted_sum[28][7:3] > 6 ? 4'd6 : weighted_sum[28][6:3]);
assign relu_out[29] = (weighted_sum[29][8]==1) ? 4'd0 : (weighted_sum[29][7:3] > 6 ? 4'd6 : weighted_sum[29][6:3]);
assign relu_out[30] = (weighted_sum[30][8]==1) ? 4'd0 : (weighted_sum[30][7:3] > 6 ? 4'd6 : weighted_sum[30][6:3]);
assign relu_out[31] = (weighted_sum[31][8]==1) ? 4'd0 : (weighted_sum[31][7:3] > 6 ? 4'd6 : weighted_sum[31][6:3]);
assign out = {relu_out[31],relu_out[30],relu_out[29],relu_out[28],relu_out[27],relu_out[26],relu_out[25],relu_out[24],relu_out[23],relu_out[22],relu_out[21],relu_out[20],relu_out[19],relu_out[18],relu_out[17],relu_out[16],relu_out[15],relu_out[14],relu_out[13],relu_out[12],relu_out[11],relu_out[10],relu_out[9],relu_out[8],relu_out[7],relu_out[6],relu_out[5],relu_out[4],relu_out[3],relu_out[2],relu_out[1],relu_out[0]};

endmodule
