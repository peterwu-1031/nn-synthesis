module fc1 (
	input [3:0] in [0:506],
	input clk,
	input rst,
	output [3:0] out [0:31]
);

logic [9:0] weighted_sum [0:31];
logic [9:0] sharing0_r, sharing0_w;
logic [9:0] sharing1_r, sharing1_w;
logic [9:0] sharing2_r, sharing2_w;
logic [9:0] sharing3_r, sharing3_w;
logic [9:0] sharing4_r, sharing4_w;
logic [9:0] sharing5_r, sharing5_w;
logic [9:0] sharing6_r, sharing6_w;
logic [9:0] sharing7_r, sharing7_w;
logic [9:0] sharing8_r, sharing8_w;
logic [9:0] sharing9_r, sharing9_w;
logic [9:0] sharing10_r, sharing10_w;
logic [9:0] sharing11_r, sharing11_w;
logic [9:0] sharing12_r, sharing12_w;
logic [9:0] sharing13_r, sharing13_w;
logic [9:0] sharing14_r, sharing14_w;
logic [9:0] sharing15_r, sharing15_w;
logic [9:0] sharing16_r, sharing16_w;
logic [9:0] sharing17_r, sharing17_w;
logic [9:0] sharing18_r, sharing18_w;
logic [9:0] sharing19_r, sharing19_w;
logic [9:0] sharing20_r, sharing20_w;
logic [9:0] sharing21_r, sharing21_w;
logic [9:0] sharing22_r, sharing22_w;
logic [9:0] sharing23_r, sharing23_w;
logic [9:0] sharing24_r, sharing24_w;
logic [9:0] sharing25_r, sharing25_w;
logic [9:0] sharing26_r, sharing26_w;
logic [9:0] sharing27_r, sharing27_w;
logic [9:0] sharing28_r, sharing28_w;
logic [9:0] sharing29_r, sharing29_w;
logic [9:0] sharing30_r, sharing30_w;
logic [9:0] sharing31_r, sharing31_w;
logic [9:0] sharing32_r, sharing32_w;
logic [9:0] sharing33_r, sharing33_w;
logic [9:0] sharing34_r, sharing34_w;
logic [9:0] sharing35_r, sharing35_w;
logic [9:0] sharing36_r, sharing36_w;
logic [9:0] sharing37_r, sharing37_w;
logic [9:0] sharing38_r, sharing38_w;
logic [9:0] sharing39_r, sharing39_w;
logic [9:0] sharing40_r, sharing40_w;
logic [9:0] sharing41_r, sharing41_w;
logic [9:0] sharing42_r, sharing42_w;
logic [9:0] sharing43_r, sharing43_w;
logic [9:0] sharing44_r, sharing44_w;
logic [9:0] sharing45_r, sharing45_w;
logic [9:0] sharing46_r, sharing46_w;
logic [9:0] sharing47_r, sharing47_w;
logic [9:0] sharing48_r, sharing48_w;
logic [9:0] sharing49_r, sharing49_w;
logic [9:0] sharing50_r, sharing50_w;
logic [9:0] sharing51_r, sharing51_w;
logic [9:0] sharing52_r, sharing52_w;
logic [9:0] sharing53_r, sharing53_w;
logic [9:0] sharing54_r, sharing54_w;
logic [9:0] sharing55_r, sharing55_w;
logic [9:0] sharing56_r, sharing56_w;
logic [9:0] sharing57_r, sharing57_w;
logic [9:0] sharing58_r, sharing58_w;
logic [9:0] sharing59_r, sharing59_w;
logic [9:0] sharing60_r, sharing60_w;
logic [9:0] sharing61_r, sharing61_w;
logic [9:0] sharing62_r, sharing62_w;
logic [9:0] sharing63_r, sharing63_w;
logic [9:0] sharing64_r, sharing64_w;
logic [9:0] sharing65_r, sharing65_w;
logic [9:0] sharing66_r, sharing66_w;
logic [9:0] sharing67_r, sharing67_w;
logic [9:0] sharing68_r, sharing68_w;
logic [9:0] sharing69_r, sharing69_w;
logic [9:0] sharing70_r, sharing70_w;
logic [9:0] sharing71_r, sharing71_w;
logic [9:0] sharing72_r, sharing72_w;
logic [9:0] sharing73_r, sharing73_w;
logic [9:0] sharing74_r, sharing74_w;
logic [9:0] sharing75_r, sharing75_w;
logic [9:0] sharing76_r, sharing76_w;
logic [9:0] sharing77_r, sharing77_w;
logic [9:0] sharing78_r, sharing78_w;
logic [9:0] sharing79_r, sharing79_w;
logic [9:0] sharing80_r, sharing80_w;
logic [9:0] sharing81_r, sharing81_w;
logic [9:0] sharing82_r, sharing82_w;
logic [9:0] sharing83_r, sharing83_w;
logic [9:0] sharing84_r, sharing84_w;
logic [9:0] sharing85_r, sharing85_w;
logic [9:0] sharing86_r, sharing86_w;
logic [9:0] sharing87_r, sharing87_w;
logic [9:0] sharing88_r, sharing88_w;
logic [9:0] sharing89_r, sharing89_w;
logic [9:0] sharing90_r, sharing90_w;
logic [9:0] sharing91_r, sharing91_w;
logic [9:0] sharing92_r, sharing92_w;
logic [9:0] sharing93_r, sharing93_w;
logic [9:0] sharing94_r, sharing94_w;
logic [9:0] sharing95_r, sharing95_w;
logic [9:0] sharing96_r, sharing96_w;
logic [9:0] sharing97_r, sharing97_w;
logic [9:0] sharing98_r, sharing98_w;
logic [9:0] sharing99_r, sharing99_w;
logic [9:0] sharing100_r, sharing100_w;
logic [9:0] sharing101_r, sharing101_w;
logic [9:0] sharing102_r, sharing102_w;
logic [9:0] sharing103_r, sharing103_w;
logic [9:0] sharing104_r, sharing104_w;
logic [9:0] sharing105_r, sharing105_w;
logic [9:0] sharing106_r, sharing106_w;
logic [9:0] sharing107_r, sharing107_w;
logic [9:0] sharing108_r, sharing108_w;
logic [9:0] sharing109_r, sharing109_w;
logic [9:0] sharing110_r, sharing110_w;
logic [9:0] sharing111_r, sharing111_w;
logic [9:0] sharing112_r, sharing112_w;
logic [9:0] sharing113_r, sharing113_w;
logic [9:0] sharing114_r, sharing114_w;
logic [9:0] sharing115_r, sharing115_w;
logic [9:0] sharing116_r, sharing116_w;
logic [9:0] sharing117_r, sharing117_w;
logic [9:0] sharing118_r, sharing118_w;
logic [9:0] sharing119_r, sharing119_w;
logic [9:0] sharing120_r, sharing120_w;
logic [9:0] sharing121_r, sharing121_w;
logic [9:0] sharing122_r, sharing122_w;
logic [9:0] sharing123_r, sharing123_w;
logic [9:0] sharing124_r, sharing124_w;
logic [9:0] sharing125_r, sharing125_w;
logic [9:0] sharing126_r, sharing126_w;
logic [9:0] sharing127_r, sharing127_w;
logic [9:0] sharing128_r, sharing128_w;
logic [9:0] sharing129_r, sharing129_w;
logic [9:0] sharing130_r, sharing130_w;
logic [9:0] sharing131_r, sharing131_w;
logic [9:0] sharing132_r, sharing132_w;
logic [9:0] sharing133_r, sharing133_w;
logic [9:0] sharing134_r, sharing134_w;
logic [9:0] sharing135_r, sharing135_w;
logic [9:0] sharing136_r, sharing136_w;
logic [9:0] sharing137_r, sharing137_w;
logic [9:0] sharing138_r, sharing138_w;
logic [9:0] sharing139_r, sharing139_w;
logic [9:0] sharing140_r, sharing140_w;
logic [9:0] sharing141_r, sharing141_w;
logic [9:0] sharing142_r, sharing142_w;
logic [9:0] sharing143_r, sharing143_w;
logic [9:0] sharing144_r, sharing144_w;
logic [9:0] sharing145_r, sharing145_w;
logic [9:0] sharing146_r, sharing146_w;
logic [9:0] sharing147_r, sharing147_w;
logic [9:0] sharing148_r, sharing148_w;
logic [9:0] sharing149_r, sharing149_w;
logic [9:0] sharing150_r, sharing150_w;
logic [9:0] sharing151_r, sharing151_w;
logic [9:0] sharing152_r, sharing152_w;
logic [9:0] sharing153_r, sharing153_w;
logic [9:0] sharing154_r, sharing154_w;
logic [9:0] sharing155_r, sharing155_w;
logic [9:0] sharing156_r, sharing156_w;
logic [9:0] sharing157_r, sharing157_w;
logic [9:0] sharing158_r, sharing158_w;
logic [9:0] sharing159_r, sharing159_w;
logic [9:0] sharing160_r, sharing160_w;
logic [9:0] sharing161_r, sharing161_w;
logic [9:0] sharing162_r, sharing162_w;
logic [9:0] sharing163_r, sharing163_w;
logic [9:0] sharing164_r, sharing164_w;
logic [9:0] sharing165_r, sharing165_w;
logic [9:0] sharing166_r, sharing166_w;
logic [9:0] sharing167_r, sharing167_w;
logic [9:0] sharing168_r, sharing168_w;
logic [9:0] sharing169_r, sharing169_w;
logic [9:0] sharing170_r, sharing170_w;
logic [9:0] sharing171_r, sharing171_w;
logic [9:0] sharing172_r, sharing172_w;
logic [9:0] sharing173_r, sharing173_w;
logic [9:0] sharing174_r, sharing174_w;
logic [9:0] sharing175_r, sharing175_w;
logic [9:0] sharing176_r, sharing176_w;
logic [9:0] sharing177_r, sharing177_w;
logic [9:0] sharing178_r, sharing178_w;
logic [9:0] sharing179_r, sharing179_w;
logic [9:0] sharing180_r, sharing180_w;
logic [9:0] sharing181_r, sharing181_w;
logic [9:0] sharing182_r, sharing182_w;
logic [9:0] sharing183_r, sharing183_w;
logic [9:0] sharing184_r, sharing184_w;
logic [9:0] sharing185_r, sharing185_w;
logic [9:0] sharing186_r, sharing186_w;
logic [9:0] sharing187_r, sharing187_w;
logic [9:0] sharing188_r, sharing188_w;
logic [9:0] sharing189_r, sharing189_w;
logic [9:0] sharing190_r, sharing190_w;
logic [9:0] sharing191_r, sharing191_w;
logic [9:0] sharing192_r, sharing192_w;
logic [9:0] sharing193_r, sharing193_w;
logic [9:0] sharing194_r, sharing194_w;
logic [9:0] sharing195_r, sharing195_w;
logic [9:0] sharing196_r, sharing196_w;
logic [9:0] sharing197_r, sharing197_w;
logic [9:0] sharing198_r, sharing198_w;
logic [9:0] sharing199_r, sharing199_w;
logic [9:0] sharing200_r, sharing200_w;
logic [9:0] sharing201_r, sharing201_w;
logic [9:0] sharing202_r, sharing202_w;
logic [9:0] sharing203_r, sharing203_w;
logic [9:0] sharing204_r, sharing204_w;
logic [9:0] sharing205_r, sharing205_w;
logic [9:0] sharing206_r, sharing206_w;
logic [9:0] sharing207_r, sharing207_w;
logic [9:0] sharing208_r, sharing208_w;
logic [9:0] sharing209_r, sharing209_w;
logic [9:0] sharing210_r, sharing210_w;
logic [9:0] sharing211_r, sharing211_w;
logic [9:0] sharing212_r, sharing212_w;
logic [9:0] sharing213_r, sharing213_w;
logic [9:0] sharing214_r, sharing214_w;
logic [9:0] sharing215_r, sharing215_w;
logic [9:0] sharing216_r, sharing216_w;
logic [9:0] sharing217_r, sharing217_w;
logic [9:0] sharing218_r, sharing218_w;
logic [9:0] sharing219_r, sharing219_w;
logic [9:0] sharing220_r, sharing220_w;
logic [9:0] sharing221_r, sharing221_w;
logic [9:0] sharing222_r, sharing222_w;
logic [9:0] sharing223_r, sharing223_w;
logic [9:0] sharing224_r, sharing224_w;
logic [9:0] sharing225_r, sharing225_w;
logic [9:0] sharing226_r, sharing226_w;
logic [9:0] sharing227_r, sharing227_w;
logic [9:0] sharing228_r, sharing228_w;
logic [9:0] sharing229_r, sharing229_w;
logic [9:0] sharing230_r, sharing230_w;
logic [9:0] sharing231_r, sharing231_w;
logic [9:0] sharing232_r, sharing232_w;
logic [9:0] sharing233_r, sharing233_w;
logic [9:0] sharing234_r, sharing234_w;
logic [9:0] sharing235_r, sharing235_w;
logic [9:0] sharing236_r, sharing236_w;
logic [9:0] sharing237_r, sharing237_w;
logic [9:0] sharing238_r, sharing238_w;
logic [9:0] sharing239_r, sharing239_w;
logic [9:0] sharing240_r, sharing240_w;
logic [9:0] sharing241_r, sharing241_w;
logic [9:0] sharing242_r, sharing242_w;
logic [9:0] sharing243_r, sharing243_w;
logic [9:0] sharing244_r, sharing244_w;
logic [9:0] sharing245_r, sharing245_w;
logic [9:0] sharing246_r, sharing246_w;
logic [9:0] sharing247_r, sharing247_w;
logic [9:0] sharing248_r, sharing248_w;
logic [9:0] sharing249_r, sharing249_w;
logic [9:0] sharing250_r, sharing250_w;
logic [9:0] sharing251_r, sharing251_w;
logic [9:0] sharing252_r, sharing252_w;
logic [9:0] sharing253_r, sharing253_w;
logic [9:0] sharing254_r, sharing254_w;
logic [9:0] sharing255_r, sharing255_w;

always_comb begin
	sharing0_w = $signed(in[128])+$signed(in[64])+$signed(in[448])+$signed(in[256])+$signed(in[417])+$signed(in[321])+$signed(in[449])+$signed(in[290])+$signed(in[322])+$signed(in[163])+$signed(in[67])+$signed(in[323])+$signed(in[318])+$signed({in[166],1'b0})+$signed(in[454])+$signed(in[70])+$signed(in[38])+$signed(in[166])+$signed(in[71])+$signed(in[167])+$signed(in[319])+$signed(in[233])+$signed({in[428],1'b0})+$signed(in[333])+$signed({in[430],1'b0})+$signed({in[334],1'b0})+$signed({in[335],1'b0})+$signed(in[207])+$signed(in[336])+$signed(in[17])+$signed({in[402],1'b0})+$signed(in[18])+$signed(in[434])+$signed(in[82])+$signed({in[243],1'b0})+$signed(in[83])+$signed(in[148])+$signed(in[213])+$signed(in[501])+$signed(in[406])+$signed(in[150])+$signed({in[503],1'b0})+$signed(in[376])+$signed(in[504])+$signed({in[153],1'b0})+$signed(in[505])+$signed(in[218])+$signed(in[94])+$signed(in[61])+$signed(in[62])+$signed({in[415],1'b0})+$signed(in[383])+$signed(-in[353])+$signed(-in[259])+$signed(-in[131])+$signed(-{in[356],1'b0})+$signed(-in[198])+$signed(-in[102])+$signed(-in[135])+$signed(-in[199])+$signed(-in[263])+$signed(-in[136])+$signed(-in[40])+$signed(-in[9])+$signed(-in[267])+$signed(-in[15])+$signed(-in[271])+$signed(-in[272])+$signed(-{in[17],2'b0})+$signed(-in[241])+$signed(-{in[18],2'b0})+$signed(-{in[19],2'b0})+$signed(-in[211])+$signed(-in[467])+$signed(-{in[23],1'b0})+$signed(-in[90])+$signed(-in[474])+$signed(-in[187])+$signed(-in[123])+$signed(-in[284])+$signed(-in[124])+$signed(-in[254])+$signed(-in[190]);
	sharing1_w = $signed(in[35])+$signed(in[132])+$signed(in[292])+$signed(in[293])+$signed(in[358])+$signed(in[456])+$signed(in[105])+$signed(in[457])+$signed(in[106])+$signed({in[492],1'b0})+$signed(in[462])+$signed(in[400])+$signed(in[469])+$signed(in[470])+$signed(in[311])+$signed(in[120])+$signed(in[440])+$signed(in[345])+$signed(in[441])+$signed(in[154])+$signed(in[314])+$signed(in[506])+$signed(in[478])+$signed(-in[129])+$signed(-in[65])+$signed(-in[225])+$signed(-in[390])+$signed(-in[103])+$signed(-in[455])+$signed(-in[327])+$signed(-in[392])+$signed(-in[41])+$signed(-in[425])+$signed(-in[44])+$signed(-in[429])+$signed(-in[238])+$signed(-in[16])+$signed(-in[276])+$signed(-in[437])+$signed(-in[22])+$signed(-in[54])+$signed(-in[438])+$signed(-in[56])+$signed(-in[88])+$signed(-in[27])+$signed(-in[381]);
	sharing2_w = $signed({in[128],1'b0})+$signed(in[64])+$signed(in[128])+$signed(in[63])+$signed(in[481])+$signed(in[129])+$signed({in[482],1'b0})+$signed(in[450])+$signed(in[354])+$signed(in[35])+$signed(in[483])+$signed({in[132],1'b0})+$signed({in[356],1'b0})+$signed({in[133],1'b0})+$signed(in[485])+$signed({in[357],1'b0})+$signed({in[454],1'b0})+$signed(in[358])+$signed(in[103])+$signed(in[487])+$signed({in[297],1'b0})+$signed(in[490])+$signed(in[427])+$signed(in[428])+$signed(in[76])+$signed(in[332])+$signed({in[77],1'b0})+$signed(in[479])+$signed(in[399])+$signed({in[368],1'b0})+$signed({in[369],1'b0})+$signed(in[17])+$signed(in[241])+$signed({in[18],1'b0})+$signed({in[466],1'b0})+$signed({in[370],1'b0})+$signed({in[19],1'b0})+$signed(in[19])+$signed(in[51])+$signed(in[307])+$signed(in[467])+$signed(in[20])+$signed({in[371],1'b0})+$signed({in[115],1'b0})+$signed({in[116],1'b0})+$signed(in[437])+$signed(in[469])+$signed({in[372],1'b0})+$signed({in[310],1'b0})+$signed({in[470],1'b0})+$signed({in[373],1'b0})+$signed(in[501])+$signed(in[246])+$signed(in[471])+$signed(in[374])+$signed(in[152])+$signed(in[440])+$signed(in[472])+$signed(in[120])+$signed(in[345])+$signed(in[121])+$signed(in[90])+$signed(in[474])+$signed(in[412])+$signed(in[413])+$signed({in[478],1'b0})+$signed(in[382])+$signed({in[127],1'b0})+$signed(in[223])+$signed(-in[256])+$signed(-in[99])+$signed(-in[101])+$signed(-in[293])+$signed(-in[262])+$signed(-in[102])+$signed(-in[390])+$signed(-in[166])+$signed(-in[391])+$signed(-in[40])+$signed(-in[41])+$signed(-in[73])+$signed(-in[78])+$signed(-in[79])+$signed(-in[432])+$signed(-in[403])+$signed(-in[275])+$signed(-in[52])+$signed(-in[85])+$signed(-in[278])+$signed(-in[86])+$signed(-in[87])+$signed(-in[27])+$signed(-in[443])+$signed(-{in[92],1'b0})+$signed(-in[317])+$signed(-{in[158],1'b0})+$signed(-in[446])+$signed(-in[95]);
	sharing3_w = $signed(in[258])+$signed(in[276])+$signed(in[377])+$signed(-in[336])+$signed(-in[389])+$signed(-in[113])+$signed(-in[401])+$signed(-in[505])+$signed(-in[107])+$signed(-in[411])+$signed(-in[108])+$signed(-in[204])+$signed(-in[324])+$signed(-in[388])+$signed(-in[189])+$signed(-in[495])+$signed(-in[167]);
	sharing4_w = $signed(in[256])+$signed(in[449])+$signed(in[193])+$signed(in[225])+$signed(in[386])+$signed(in[450])+$signed(in[99])+$signed(in[291])+$signed(in[483])+$signed(in[36])+$signed(in[229])+$signed(in[69])+$signed(in[166])+$signed(in[423])+$signed(in[167])+$signed(in[199])+$signed(in[447])+$signed(in[205])+$signed(in[77])+$signed(in[269])+$signed(in[206])+$signed(in[238])+$signed(in[432])+$signed(in[81])+$signed({in[436],1'b0})+$signed(in[212])+$signed(in[214])+$signed(in[22])+$signed(in[438])+$signed(in[279])+$signed(in[375])+$signed(in[217])+$signed(in[282])+$signed(in[411])+$signed(in[412])+$signed(in[317])+$signed(in[446])+$signed(in[415])+$signed(-in[344])+$signed(-in[440])+$signed(-in[441])+$signed(-in[473])+$signed(-in[17])+$signed(-in[58])+$signed(-in[491])+$signed(-in[356])+$signed(-in[357])+$signed(-in[6])+$signed(-in[7]);
	sharing5_w = $signed(in[224])+$signed(in[417])+$signed(in[258])+$signed(in[419])+$signed(in[131])+$signed(in[68])+$signed(in[134])+$signed(in[454])+$signed(in[422])+$signed(in[359])+$signed(in[40])+$signed(in[232])+$signed(in[392])+$signed(in[42])+$signed(in[43])+$signed({in[76],1'b0})+$signed(in[332])+$signed(in[79])+$signed(in[399])+$signed(in[463])+$signed(in[304])+$signed(in[371])+$signed(in[467])+$signed({in[404],1'b0})+$signed(in[116])+$signed(in[244])+$signed(in[500])+$signed(in[53])+$signed(in[245])+$signed(in[373])+$signed({in[54],1'b0})+$signed(in[405])+$signed(in[406])+$signed(in[469])+$signed(in[501])+$signed(in[56])+$signed(in[472])+$signed(in[121])+$signed(in[345])+$signed(in[30])+$signed(in[27])+$signed({in[60],1'b0})+$signed(in[380])+$signed({in[61],1'b0})+$signed({in[413],1'b0})+$signed({in[414],1'b0})+$signed(in[62])+$signed({in[63],1'b0})+$signed(in[383])+$signed(-in[24])+$signed(-in[264])+$signed(-in[448])+$signed(-in[288])+$signed(-in[280])+$signed(-in[153])+$signed(-in[506])+$signed(-in[107])+$signed(-in[187])+$signed(-in[268])+$signed(-in[84])+$signed(-in[252])+$signed(-in[284])+$signed(-in[479])+$signed(-in[191])+$signed(-in[503])+$signed(-in[190])+$signed(-in[335]);
	sharing6_w = $signed(in[416])+$signed(in[164])+$signed(in[165])+$signed({in[166],1'b0})+$signed(in[70])+$signed(in[422])+$signed({in[423],1'b0})+$signed(in[40])+$signed(in[72])+$signed(in[200])+$signed(in[424])+$signed(in[201])+$signed(in[265])+$signed(in[297])+$signed(in[457])+$signed(in[459])+$signed(in[415])+$signed(in[460])+$signed(in[237])+$signed(in[239])+$signed(in[367])+$signed(in[399])+$signed(in[431])+$signed(in[112])+$signed(in[495])+$signed(in[17])+$signed(in[113])+$signed(in[241])+$signed(in[401])+$signed(in[18])+$signed(in[115])+$signed(in[403])+$signed(in[376])+$signed(in[441])+$signed(in[410])+$signed({in[251],1'b0})+$signed(in[59])+$signed(in[411])+$signed(in[443])+$signed(in[252])+$signed(in[413])+$signed(in[30])+$signed(in[127])+$signed(-in[153])+$signed(-in[217])+$signed(-in[89])+$signed(-in[426])+$signed(-in[490])+$signed(-in[50])+$signed(-in[323])+$signed(-in[491])+$signed(-in[147])+$signed(-in[219])+$signed(-in[492])+$signed(-in[468])+$signed(-in[220])+$signed(-in[477])+$signed(-in[358])+$signed(-in[7])+$signed(-in[135]);
	sharing7_w = $signed(in[385])+$signed(in[449])+$signed(in[35])+$signed(in[483])+$signed(in[68])+$signed(in[484])+$signed(in[485])+$signed(in[39])+$signed(in[391])+$signed(in[303])+$signed(in[368])+$signed(in[369])+$signed(in[466])+$signed(in[467])+$signed(in[405])+$signed(in[53])+$signed(in[407])+$signed(in[280])+$signed(in[408])+$signed(in[379])+$signed(in[380])+$signed(-in[192])+$signed(-in[320])+$signed(-in[193])+$signed(-in[353])+$signed(-in[354])+$signed(-in[355])+$signed(-in[356])+$signed(-in[6])+$signed(-in[198])+$signed(-in[136])+$signed(-in[360])+$signed(-in[456])+$signed(-in[9])+$signed(-in[138])+$signed(-in[206])+$signed(-in[270])+$signed(-in[15])+$signed(-in[432])+$signed(-in[83])+$signed(-in[149])+$signed(-in[469])+$signed(-in[150])+$signed(-in[470])+$signed(-in[502])+$signed(-{in[23],1'b0})+$signed(-in[471])+$signed(-in[216])+$signed(-in[186])+$signed(-in[187])+$signed(-in[475])+$signed(-in[28])+$signed(-in[189])+$signed(-in[190]);
	sharing8_w = $signed(in[192])+$signed(in[193])+$signed(in[353])+$signed(in[450])+$signed(in[100])+$signed(in[357])+$signed(in[389])+$signed(in[382])+$signed({in[102],1'b0})+$signed({in[454],1'b0})+$signed({in[199],1'b0})+$signed(in[423])+$signed(in[487])+$signed(in[488])+$signed({in[393],1'b0})+$signed(in[9])+$signed(in[41])+$signed(in[266])+$signed(in[269])+$signed(in[270])+$signed(in[398])+$signed(in[271])+$signed(in[399])+$signed({in[272],1'b0})+$signed(in[368])+$signed(in[369])+$signed({in[18],1'b0})+$signed(in[370])+$signed(in[402])+$signed(in[19])+$signed(in[115])+$signed(in[371])+$signed(in[403])+$signed(in[372])+$signed(in[277])+$signed(in[437])+$signed({in[22],1'b0})+$signed({in[374],1'b0})+$signed(in[406])+$signed(in[438])+$signed({in[23],1'b0})+$signed(in[439])+$signed(in[24])+$signed(in[281])+$signed(in[187])+$signed(in[253])+$signed(in[189])+$signed(in[318])+$signed(in[191])+$signed(-in[152])+$signed(-in[105])+$signed(-in[457])+$signed(-in[505])+$signed(-in[481])+$signed(-in[154])+$signed(-in[302])+$signed(-in[419])+$signed(-in[323])+$signed(-in[491])+$signed(-in[324])+$signed(-in[140])+$signed(-in[492])+$signed(-{in[165],1'b0})+$signed(-{in[421],1'b0})+$signed(-in[334])+$signed(-in[430])+$signed(-in[167]);
	sharing9_w = $signed({in[161],1'b0})+$signed(in[129])+$signed(in[162])+$signed(in[387])+$signed(in[132])+$signed(in[484])+$signed(in[5])+$signed(in[7])+$signed(in[327])+$signed(in[296])+$signed(in[328])+$signed(in[329])+$signed(in[361])+$signed(in[362])+$signed(in[43])+$signed(in[331])+$signed(in[236])+$signed(in[493])+$signed(in[238])+$signed(in[304])+$signed(in[400])+$signed(in[49])+$signed(in[497])+$signed(in[146])+$signed(in[119])+$signed(in[407])+$signed(in[120])+$signed(in[344])+$signed(in[57])+$signed(in[249])+$signed(in[58])+$signed(in[314])+$signed(in[411])+$signed(in[478])+$signed(in[127])+$signed(-in[288])+$signed(-in[97])+$signed(-in[225])+$signed(-in[66])+$signed(-in[37])+$signed(-in[166])+$signed(-in[458])+$signed(-in[141])+$signed(-in[206])+$signed(-in[462])+$signed(-in[111])+$signed(-in[432])+$signed(-in[401])+$signed(-in[433])+$signed(-in[82])+$signed(-in[242])+$signed(-in[434])+$signed(-in[218])+$signed(-in[220])+$signed(-in[444])+$signed(-in[93])+$signed(-in[255]);
	sharing10_w = $signed(in[32])+$signed(in[224])+$signed({in[449],1'b0})+$signed(in[289])+$signed(in[257])+$signed(in[321])+$signed(in[34])+$signed({in[451],1'b0})+$signed(in[131])+$signed(in[35])+$signed(in[99])+$signed({in[452],1'b0})+$signed(in[36])+$signed(in[356])+$signed(in[357])+$signed(in[358])+$signed(in[393])+$signed(in[394])+$signed(in[138])+$signed(in[330])+$signed({in[43],1'b0})+$signed(in[108])+$signed(in[492])+$signed(in[269])+$signed(in[141])+$signed(in[237])+$signed(in[334])+$signed({in[368],1'b0})+$signed({in[466],1'b0})+$signed(in[18])+$signed(in[370])+$signed(in[51])+$signed(in[115])+$signed(in[371])+$signed({in[212],1'b0})+$signed(in[276])+$signed(in[308])+$signed(in[116])+$signed({in[437],1'b0})+$signed(in[405])+$signed(in[309])+$signed(in[29])+$signed({in[438],1'b0})+$signed(in[310])+$signed({in[374],1'b0})+$signed(in[502])+$signed({in[439],1'b0})+$signed(in[407])+$signed(in[215])+$signed(in[408])+$signed(in[504])+$signed({in[30],1'b0})+$signed(in[250])+$signed(in[285])+$signed({in[478],1'b0})+$signed(in[446])+$signed(in[383])+$signed(-in[64])+$signed(-in[416])+$signed(-{in[65],1'b0})+$signed(-in[388])+$signed(-in[390])+$signed(-in[327])+$signed(-in[71])+$signed(-in[265])+$signed(-in[458])+$signed(-in[106])+$signed(-in[75])+$signed(-in[76])+$signed(-in[429])+$signed(-in[78])+$signed(-in[16])+$signed(-in[400])+$signed(-in[496])+$signed(-in[401])+$signed(-in[403])+$signed(-in[52])+$signed(-in[246])+$signed(-in[61])+$signed(-in[411])+$signed(-in[59])+$signed(-in[315])+$signed(-in[60])+$signed(-in[413])+$signed(-in[414])+$signed(-{in[415],1'b0})+$signed(-in[63]);
	sharing11_w = $signed(in[264])+$signed(in[314])+$signed(in[38])+$signed(in[302])+$signed(in[54])+$signed(in[427])+$signed(in[292])+$signed(in[460])+$signed(in[404])+$signed(in[158])+$signed(in[391])+$signed(-in[456])+$signed(-in[424])+$signed(-in[345])+$signed(-in[457])+$signed(-in[119])+$signed(-in[282])+$signed(-in[469])+$signed(-in[387])+$signed(-in[163])+$signed(-in[107])+$signed(-in[83])+$signed(-in[253])+$signed(-in[278])+$signed(-in[471]);
	sharing12_w = $signed(in[288])+$signed(in[417])+$signed(in[226])+$signed(in[290])+$signed(in[484])+$signed(in[262])+$signed(in[135])+$signed(in[231])+$signed({in[264],1'b0})+$signed(in[490])+$signed(in[140])+$signed(in[268])+$signed(in[237])+$signed(in[141])+$signed(in[301])+$signed(in[78])+$signed(in[142])+$signed(in[145])+$signed(in[241])+$signed(in[305])+$signed(in[434])+$signed(in[243])+$signed(in[435])+$signed(in[276])+$signed(in[279])+$signed(in[249])+$signed(in[317])+$signed({in[250],1'b0})+$signed({in[251],1'b0})+$signed(in[315])+$signed({in[252],1'b0})+$signed(in[316])+$signed(in[477])+$signed(in[158])+$signed(in[255])+$signed(-in[481])+$signed(-in[450])+$signed(-in[388])+$signed(-in[414])+$signed(-in[455])+$signed(-in[456])+$signed(-in[105])+$signed(-in[425])+$signed(-in[426])+$signed(-in[460])+$signed(-in[367])+$signed(-in[368])+$signed(-{in[434],2'b0})+$signed(-in[83])+$signed(-{in[436],1'b0})+$signed(-in[85])+$signed(-in[438])+$signed(-in[119])+$signed(-in[439])+$signed(-in[220])+$signed(-in[30]);
	sharing13_w = $signed(in[258])+$signed(in[291])+$signed(in[387])+$signed(in[36])+$signed(in[229])+$signed(in[37])+$signed(in[166])+$signed(in[205])+$signed(in[270])+$signed(in[430])+$signed(in[47])+$signed(in[271])+$signed(in[431])+$signed(in[336])+$signed(in[400])+$signed(in[433])+$signed(in[503])+$signed(in[504])+$signed(in[24])+$signed(in[88])+$signed(in[216])+$signed({in[89],1'b0})+$signed(in[473])+$signed(in[505])+$signed(in[218])+$signed(in[219])+$signed({in[445],1'b0})+$signed(in[94])+$signed(in[191])+$signed(-in[97])+$signed(-in[163])+$signed(-in[67])+$signed(-in[69])+$signed(-in[70])+$signed(-in[391])+$signed(-in[394])+$signed(-in[403])+$signed(-in[467])+$signed(-in[116])+$signed(-in[405])+$signed(-{in[406],1'b0})+$signed(-in[86])+$signed(-in[374])+$signed(-{in[407],1'b0})+$signed(-in[440])+$signed(-{in[441],1'b0})+$signed(-in[57])+$signed(-in[410]);
	sharing14_w = $signed(in[163])+$signed(in[451])+$signed({in[422],1'b0})+$signed(in[422])+$signed(in[200])+$signed(in[264])+$signed({in[431],1'b0})+$signed(in[431])+$signed(in[463])+$signed({in[432],1'b0})+$signed(in[81])+$signed({in[82],1'b0})+$signed(in[83])+$signed(in[215])+$signed({in[408],1'b0})+$signed(in[216])+$signed(in[440])+$signed(in[57])+$signed(in[409])+$signed(in[58])+$signed(in[59])+$signed(in[379])+$signed(in[92])+$signed(in[254])+$signed(-{in[443],1'b0})+$signed(-in[95]);
	sharing15_w = $signed(in[160])+$signed(in[130])+$signed(in[356])+$signed(in[357])+$signed({in[358],1'b0})+$signed({in[454],1'b0})+$signed(in[230])+$signed(in[327])+$signed(in[455])+$signed(in[359])+$signed(in[8])+$signed(in[395])+$signed(in[492])+$signed(in[141])+$signed(in[366])+$signed(in[367])+$signed(in[48])+$signed(in[145])+$signed(in[18])+$signed({in[467],1'b0})+$signed(in[52])+$signed(in[405])+$signed(in[406])+$signed(in[119])+$signed(in[345])+$signed(in[90])+$signed(in[314])+$signed(in[30])+$signed(in[315])+$signed(in[316])+$signed(in[157])+$signed(in[158])+$signed(in[479])+$signed(-{in[64],1'b0})+$signed(-in[193])+$signed(-in[387])+$signed(-{in[421],2'b0})+$signed(-in[165])+$signed(-in[38])+$signed(-in[262])+$signed(-in[166])+$signed(-{in[71],2'b0})+$signed(-in[296])+$signed(-in[297])+$signed(-in[361])+$signed(-in[206])+$signed(-in[207])+$signed(-{in[80],2'b0})+$signed(-in[400])+$signed(-{in[51],1'b0})+$signed(-in[307])+$signed(-in[436])+$signed(-in[246])+$signed(-in[374])+$signed(-{in[375],1'b0})+$signed(-in[249])+$signed(-in[250])+$signed(-{in[252],2'b0})+$signed(-in[188])+$signed(-in[220])+$signed(-in[412])+$signed(-in[414])+$signed(-in[127]);
	sharing16_w = $signed(in[384])+$signed(in[128])+$signed(in[256])+$signed({in[225],1'b0})+$signed(in[161])+$signed(in[481])+$signed({in[258],1'b0})+$signed(in[226])+$signed(in[258])+$signed(in[451])+$signed(in[324])+$signed(in[452])+$signed({in[165],1'b0})+$signed(in[327])+$signed(in[328])+$signed(in[424])+$signed(in[425])+$signed(in[75])+$signed(in[268])+$signed({in[237],1'b0})+$signed(in[109])+$signed(in[269])+$signed(in[270])+$signed(in[334])+$signed(in[336])+$signed(in[496])+$signed(in[211])+$signed(in[403])+$signed(in[244])+$signed(in[276])+$signed(in[468])+$signed(in[213])+$signed(in[53])+$signed(in[86])+$signed(in[87])+$signed(in[279])+$signed({in[88],1'b0})+$signed(in[440])+$signed(in[89])+$signed(in[281])+$signed(in[313])+$signed(in[154])+$signed(in[442])+$signed(in[506])+$signed(in[155])+$signed({in[380],1'b0})+$signed(in[381])+$signed(in[383])+$signed(-{in[64],1'b0})+$signed(-in[344])+$signed(-in[400])+$signed(-in[389])+$signed(-in[457])+$signed(-in[361])+$signed(-in[410])+$signed(-{in[204],1'b0})+$signed(-in[4])+$signed(-in[20])+$signed(-in[493])+$signed(-in[374]);
	sharing17_w = $signed(in[8])+$signed(in[57])+$signed(in[473])+$signed(in[233])+$signed(in[202])+$signed(in[58])+$signed(in[363])+$signed(in[427])+$signed(in[219])+$signed(in[36])+$signed(in[44])+$signed(in[220])+$signed(in[5])+$signed(in[37])+$signed(in[45])+$signed(in[398])+$signed(in[63])+$signed(-in[288])+$signed(-in[416])+$signed(-in[66])+$signed(-in[259])+$signed(-in[419])+$signed(-in[229])+$signed(-in[223])+$signed(-{in[390],1'b0})+$signed(-in[454])+$signed(-in[200])+$signed(-in[43])+$signed(-in[107])+$signed(-in[76])+$signed(-in[428])+$signed(-in[301])+$signed(-in[462])+$signed(-in[431])+$signed(-in[463])+$signed(-in[79])+$signed(-{in[369],1'b0})+$signed(-in[81])+$signed(-{in[370],1'b0})+$signed(-in[434])+$signed(-in[275])+$signed(-{in[404],1'b0})+$signed(-in[52])+$signed(-in[116])+$signed(-in[277])+$signed(-{in[54],1'b0})+$signed(-in[406])+$signed(-in[55])+$signed(-in[23])+$signed(-in[407])+$signed(-in[90])+$signed(-in[378])+$signed(-{in[29],1'b0})+$signed(-in[94])+$signed(-in[31]);
	sharing18_w = $signed(in[222])+$signed(in[449])+$signed(in[129])+$signed(in[481])+$signed(in[130])+$signed(in[482])+$signed(in[445])+$signed({in[131],1'b0})+$signed(in[388])+$signed(in[327])+$signed(in[168])+$signed(in[41])+$signed(in[329])+$signed(in[425])+$signed(in[457])+$signed(in[427])+$signed(in[365])+$signed(in[238])+$signed({in[495],1'b0})+$signed(in[303])+$signed(in[207])+$signed(in[144])+$signed(in[304])+$signed(in[369])+$signed(in[497])+$signed({in[51],1'b0})+$signed(in[147])+$signed(in[148])+$signed(in[468])+$signed({in[469],1'b0})+$signed(in[375])+$signed(in[120])+$signed(in[473])+$signed(in[218])+$signed(in[314])+$signed(in[442])+$signed(in[379])+$signed(in[220])+$signed(in[253])+$signed(in[380])+$signed(in[317])+$signed({in[158],1'b0})+$signed(in[126])+$signed({in[415],1'b0})+$signed(in[95])+$signed(-in[416])+$signed(-in[65])+$signed(-in[354])+$signed(-{in[292],2'b0})+$signed(-in[165])+$signed(-in[255])+$signed(-in[103])+$signed(-in[74])+$signed(-in[202])+$signed(-{in[107],1'b0})+$signed(-in[111])+$signed(-in[271])+$signed(-in[16])+$signed(-in[464])+$signed(-in[242])+$signed(-in[243])+$signed(-in[275])+$signed(-in[244])+$signed(-in[23])+$signed(-in[24])+$signed(-in[248])+$signed(-in[506])+$signed(-in[188])+$signed(-in[412])+$signed(-in[189])+$signed(-in[414])+$signed(-in[190]);
	sharing19_w = $signed(in[357])+$signed(in[454])+$signed(in[456])+$signed(in[200])+$signed(in[33])+$signed(in[17])+$signed(in[278])+$signed({in[443],1'b0})+$signed(in[419])+$signed(in[19])+$signed(in[356])+$signed(in[420])+$signed(in[366])+$signed(in[20])+$signed(in[421])+$signed(in[276])+$signed(in[277])+$signed(in[270])+$signed(-in[206])+$signed(-in[440])+$signed(-in[97])+$signed(-in[265])+$signed(-in[266])+$signed(-in[439])+$signed(-in[164])+$signed(-in[404])+$signed(-in[53])+$signed(-in[406])+$signed(-in[462])+$signed(-in[93])+$signed(-in[191]);
	sharing20_w = $signed(in[384])+$signed(in[64])+$signed(in[192])+$signed({in[385],1'b0})+$signed(in[353])+$signed({in[386],2'b0})+$signed(in[34])+$signed(in[258])+$signed({in[387],1'b0})+$signed(in[355])+$signed(in[389])+$signed(in[358])+$signed(in[486])+$signed(in[263])+$signed(in[264])+$signed(in[424])+$signed(in[361])+$signed(in[331])+$signed(in[76])+$signed(in[397])+$signed({in[398],1'b0})+$signed({in[399],1'b0})+$signed(in[400])+$signed(in[496])+$signed(in[402])+$signed(in[19])+$signed(in[51])+$signed(in[371])+$signed({in[372],1'b0})+$signed(in[245])+$signed(in[22])+$signed(in[278])+$signed(in[374])+$signed(in[470])+$signed(in[215])+$signed(in[24])+$signed(in[472])+$signed(in[89])+$signed(in[345])+$signed(in[219])+$signed(in[475])+$signed(in[415])+$signed(-in[117])+$signed(-in[104])+$signed(-{in[41],1'b0})+$signed(-in[367])+$signed(-in[211])+$signed(-in[468])+$signed(-in[28])+$signed(-in[92])+$signed(-in[223])+$signed(-in[381])+$signed(-in[430])+$signed(-in[455]);
	sharing21_w = $signed(in[288])+$signed(in[226])+$signed(in[227])+$signed({in[388],1'b0})+$signed(in[36])+$signed(in[38])+$signed({in[232],1'b0})+$signed(in[200])+$signed(in[392])+$signed({in[233],1'b0})+$signed(in[201])+$signed(in[297])+$signed(in[393])+$signed({in[205],1'b0})+$signed(in[77])+$signed(in[302])+$signed(in[207])+$signed(in[401])+$signed(in[214])+$signed(in[61])+$signed(in[376])+$signed(in[189])+$signed(in[93])+$signed(in[62])+$signed(in[63])+$signed(-in[32])+$signed(-in[160])+$signed(-in[416])+$signed(-in[417])+$signed(-in[418])+$signed(-in[67])+$signed(-{in[229],1'b0})+$signed(-in[165])+$signed(-in[453])+$signed(-in[103])+$signed(-in[72])+$signed(-in[328])+$signed(-in[236])+$signed(-in[268])+$signed(-in[335])+$signed(-in[272])+$signed(-{in[249],1'b0})+$signed(-in[154])+$signed(-in[250])+$signed(-in[506])+$signed(-{in[59],1'b0})+$signed(-in[155])+$signed(-in[382])+$signed(-{in[159],1'b0});
	sharing22_w = $signed(in[64])+$signed(in[96])+$signed(in[225])+$signed(in[481])+$signed(in[413])+$signed({in[482],1'b0})+$signed(in[387])+$signed(in[483])+$signed(in[132])+$signed(in[388])+$signed(in[484])+$signed(in[133])+$signed(in[134])+$signed(in[423])+$signed(in[296])+$signed(in[329])+$signed(in[330])+$signed(in[331])+$signed(in[428])+$signed({in[144],1'b0})+$signed(in[400])+$signed(in[145])+$signed(in[498])+$signed(in[51])+$signed(in[84])+$signed(in[436])+$signed(in[437])+$signed(in[470])+$signed(in[471])+$signed(in[472])+$signed(in[121])+$signed(in[253])+$signed(in[254])+$signed({in[415],1'b0})+$signed(in[127])+$signed(-{in[129],1'b0})+$signed(-in[258])+$signed(-in[259])+$signed(-in[357])+$signed(-in[102])+$signed(-in[390])+$signed(-in[103])+$signed(-in[200])+$signed(-in[235])+$signed(-in[461])+$signed(-in[78])+$signed(-in[110])+$signed(-in[79])+$signed(-in[431])+$signed(-{in[304],1'b0})+$signed(-in[80])+$signed(-in[17])+$signed(-{in[466],2'b0})+$signed(-{in[116],1'b0})+$signed(-in[52])+$signed(-in[88])+$signed(-in[248])+$signed(-in[249])+$signed(-in[441])+$signed(-in[90])+$signed(-in[188])+$signed(-in[189])+$signed(-{in[479],1'b0});
	sharing23_w = $signed(in[98])+$signed(in[292])+$signed(in[263])+$signed(in[106])+$signed(in[107])+$signed(in[267])+$signed(in[366])+$signed(in[430])+$signed(in[432])+$signed(in[433])+$signed(in[467])+$signed(in[85])+$signed(in[376])+$signed(in[89])+$signed(in[314])+$signed(in[27])+$signed(in[315])+$signed(in[28])+$signed(in[284])+$signed(in[29])+$signed(-in[128])+$signed(-in[360])+$signed(-in[361])+$signed(-in[425])+$signed(-in[337])+$signed(-in[165])+$signed(-in[205])+$signed(-in[407])+$signed(-in[211])+$signed(-in[219])+$signed(-in[245])+$signed(-in[244])+$signed(-in[141])+$signed(-in[374])+$signed(-in[279])+$signed(-in[63]);
	sharing24_w = $signed(in[161])+$signed({in[388],1'b0})+$signed(in[388])+$signed(in[421])+$signed(in[389])+$signed(in[263])+$signed(in[383])+$signed({in[395],1'b0})+$signed(in[491])+$signed({in[428],1'b0})+$signed(in[44])+$signed(in[141])+$signed(in[433])+$signed(in[242])+$signed(in[275])+$signed(in[372])+$signed(in[375])+$signed(in[408])+$signed(in[315])+$signed(in[475])+$signed(in[382])+$signed(in[159])+$signed(-in[109])+$signed(-in[336])+$signed(-in[440])+$signed(-in[249])+$signed(-in[505])+$signed(-in[257])+$signed(-{in[250],2'b0})+$signed(-in[258])+$signed(-in[354])+$signed(-{in[251],1'b0})+$signed(-{in[188],1'b0})+$signed(-in[277]);
	sharing25_w = $signed(in[193])+$signed(in[386])+$signed(in[165])+$signed(in[38])+$signed(in[7])+$signed(in[167])+$signed(in[266])+$signed(in[267])+$signed(in[268])+$signed(in[205])+$signed(in[493])+$signed(in[206])+$signed(in[334])+$signed(in[399])+$signed(in[271])+$signed({in[400],1'b0})+$signed({in[401],2'b0})+$signed(in[50])+$signed({in[51],1'b0})+$signed(in[374])+$signed(in[55])+$signed(in[151])+$signed(in[439])+$signed(in[503])+$signed(in[376])+$signed({in[409],1'b0})+$signed({in[414],1'b0})+$signed(in[190])+$signed({in[415],1'b0})+$signed(in[63])+$signed(-in[224])+$signed(-in[381])+$signed(-in[129])+$signed(-in[130])+$signed(-{in[356],1'b0})+$signed(-in[223])+$signed(-{in[358],1'b0})+$signed(-{in[391],1'b0})+$signed(-in[40])+$signed(-in[456])+$signed(-in[478])+$signed(-in[297])+$signed(-in[106])+$signed(-in[362])+$signed(-in[301])+$signed(-in[366])+$signed(-{in[368],1'b0})+$signed(-{in[19],1'b0})+$signed(-in[244])+$signed(-in[468])+$signed(-{in[53],1'b0})+$signed(-in[21])+$signed(-in[54])+$signed(-in[313])+$signed(-in[345])+$signed(-in[441])+$signed(-in[506])+$signed(-in[379])+$signed(-in[443])+$signed(-{in[92],1'b0})+$signed(-in[28])+$signed(-in[380])+$signed(-in[444])+$signed(-{in[93],1'b0})+$signed(-in[29])+$signed(-in[30])+$signed(-in[31]);
	sharing26_w = $signed(in[288])+$signed(in[480])+$signed({in[129],1'b0})+$signed(in[289])+$signed(in[385])+$signed(in[130])+$signed(in[386])+$signed(in[131])+$signed(in[355])+$signed(in[453])+$signed({in[358],1'b0})+$signed({in[454],1'b0})+$signed(in[359])+$signed(in[265])+$signed(in[107])+$signed(in[447])+$signed({in[301],1'b0})+$signed(in[109])+$signed(in[302])+$signed(in[303])+$signed(in[399])+$signed(in[80])+$signed(in[51])+$signed(in[467])+$signed({in[116],1'b0})+$signed(in[372])+$signed(in[277])+$signed(in[373])+$signed(in[278])+$signed(in[310])+$signed(in[345])+$signed(in[409])+$signed(in[314])+$signed(in[411])+$signed(in[445])+$signed(in[126])+$signed(in[31])+$signed(-{in[192],1'b0})+$signed(-in[416])+$signed(-in[481])+$signed(-in[66])+$signed(-in[68])+$signed(-in[197])+$signed(-in[6])+$signed(-in[327])+$signed(-in[71])+$signed(-in[9])+$signed(-in[41])+$signed(-in[203])+$signed(-in[429])+$signed(-{in[495],1'b0})+$signed(-in[241])+$signed(-in[403])+$signed(-in[404])+$signed(-in[85])+$signed(-in[53])+$signed(-in[54])+$signed(-in[55])+$signed(-in[23])+$signed(-in[24])+$signed(-in[89])+$signed(-in[28])+$signed(-in[188])+$signed(-{in[190],1'b0})+$signed(-in[254])+$signed(-in[255]);
	sharing27_w = $signed(in[320])+$signed(in[387])+$signed(in[36])+$signed({in[37],1'b0})+$signed({in[165],1'b0})+$signed({in[166],1'b0})+$signed(in[391])+$signed(in[489])+$signed(in[426])+$signed(in[430])+$signed(in[431])+$signed(in[207])+$signed({in[336],1'b0})+$signed(in[308])+$signed(in[438])+$signed({in[503],1'b0})+$signed(in[504])+$signed({in[505],1'b0})+$signed(in[153])+$signed(in[249])+$signed(in[154])+$signed(in[155])+$signed({in[252],1'b0})+$signed(-in[160])+$signed(-in[63])+$signed(-in[290])+$signed(-in[418])+$signed(-in[452])+$signed(-in[199])+$signed(-in[200])+$signed(-in[330])+$signed(-in[428])+$signed(-in[111])+$signed(-in[15])+$signed(-in[497])+$signed(-in[498])+$signed(-in[83])+$signed(-in[435])+$signed(-in[499])+$signed(-in[246])+$signed(-in[408])+$signed(-in[440])+$signed(-in[157])+$signed(-in[414])+$signed(-{in[415],1'b0})+$signed(-in[159]);
	sharing28_w = $signed(in[64])+$signed(in[448])+$signed(in[449])+$signed(in[450])+$signed(in[98])+$signed(in[355])+$signed(in[4])+$signed({in[255],1'b0})+$signed(in[229])+$signed(in[37])+$signed(in[223])+$signed(in[423])+$signed(in[202])+$signed({in[267],1'b0})+$signed(in[267])+$signed({in[205],1'b0})+$signed(in[461])+$signed(in[304])+$signed(in[464])+$signed(in[84])+$signed(in[116])+$signed(in[212])+$signed({in[85],1'b0})+$signed({in[23],1'b0})+$signed(in[23])+$signed(in[407])+$signed({in[24],1'b0})+$signed({in[280],1'b0})+$signed(in[408])+$signed(in[473])+$signed(in[122])+$signed(in[218])+$signed({in[187],1'b0})+$signed(in[475])+$signed(in[92])+$signed(in[188])+$signed({in[254],1'b0})+$signed({in[191],1'b0})+$signed(in[191])+$signed(-in[272])+$signed(-in[416])+$signed(-in[345])+$signed(-in[82])+$signed(-in[75])+$signed(-in[259])+$signed(-in[235])+$signed(-in[275])+$signed(-in[411])+$signed(-in[60])+$signed(-in[62])+$signed(-in[165])+$signed(-in[390])+$signed(-in[239])+$signed(-in[30])+$signed(-in[271]);
	sharing29_w = $signed(in[160])+$signed(in[161])+$signed(in[481])+$signed(in[413])+$signed(in[66])+$signed(in[34])+$signed(in[162])+$signed(in[354])+$signed(in[35])+$signed(in[71])+$signed(in[455])+$signed(in[391])+$signed(in[104])+$signed(in[296])+$signed(in[328])+$signed(in[73])+$signed(in[297])+$signed(in[329])+$signed(in[425])+$signed(in[249])+$signed(in[285])+$signed(in[158])+$signed(-in[96])+$signed(-in[324])+$signed(-in[292])+$signed(-{in[389],1'b0})+$signed(-in[453])+$signed(-in[293])+$signed(-{in[454],1'b0})+$signed(-{in[492],1'b0})+$signed(-in[428])+$signed(-in[335])+$signed(-in[112])+$signed(-in[336])+$signed(-in[337])+$signed(-in[401])+$signed(-in[465])+$signed(-in[50])+$signed(-in[402])+$signed(-in[434])+$signed(-{in[505],1'b0})+$signed(-in[281])+$signed(-in[506])+$signed(-in[155])+$signed(-in[414]);
	sharing30_w = $signed(in[256])+$signed(in[224])+$signed(in[481])+$signed(in[257])+$signed(in[132])+$signed({in[454],1'b0})+$signed(in[358])+$signed({in[391],1'b0})+$signed(in[327])+$signed(in[455])+$signed(in[392])+$signed(in[40])+$signed(in[232])+$signed(in[393])+$signed(in[41])+$signed(in[457])+$signed(in[266])+$signed(in[462])+$signed(in[366])+$signed(in[112])+$signed(in[496])+$signed(in[369])+$signed(in[242])+$signed({in[243],1'b0})+$signed(in[275])+$signed(in[435])+$signed(in[467])+$signed({in[244],1'b0})+$signed(in[276])+$signed(in[468])+$signed({in[245],1'b0})+$signed(in[118])+$signed(in[375])+$signed({in[378],1'b0})+$signed(in[442])+$signed(in[315])+$signed(in[443])+$signed(in[379])+$signed(in[124])+$signed({in[61],1'b0})+$signed(in[223])+$signed(-{in[192],1'b0})+$signed(-in[353])+$signed(-in[386])+$signed(-in[354])+$signed(-in[259])+$signed(-in[227])+$signed(-{in[388],2'b0})+$signed(-in[4])+$signed(-in[36])+$signed(-in[164])+$signed(-in[324])+$signed(-in[5])+$signed(-in[69])+$signed(-in[6])+$signed(-in[167])+$signed(-in[200])+$signed(-in[360])+$signed(-in[9])+$signed(-in[201])+$signed(-in[361])+$signed(-in[10])+$signed(-in[298])+$signed(-in[202])+$signed(-in[362])+$signed(-in[203])+$signed(-in[141])+$signed(-in[205])+$signed(-in[206])+$signed(-in[15])+$signed(-in[207])+$signed(-in[16])+$signed(-in[81])+$signed(-in[18])+$signed(-in[213])+$signed(-in[373])+$signed(-in[342])+$signed(-in[374])+$signed(-{in[375],2'b0})+$signed(-{in[23],1'b0})+$signed(-in[311])+$signed(-in[343])+$signed(-in[186])+$signed(-{in[187],1'b0})+$signed(-{in[188],1'b0})+$signed(-{in[189],1'b0})+$signed(-in[285])+$signed(-{in[190],1'b0})+$signed(-{in[191],1'b0})+$signed(-in[31]);
	sharing31_w = $signed(in[384])+$signed(in[417])+$signed(in[226])+$signed(in[67])+$signed(in[100])+$signed(in[197])+$signed(in[101])+$signed(in[414])+$signed(in[263])+$signed(in[295])+$signed(in[427])+$signed(in[459])+$signed(in[301])+$signed(in[270])+$signed(in[430])+$signed(in[79])+$signed(in[271])+$signed(in[239])+$signed(in[80])+$signed(in[400])+$signed(in[52])+$signed(in[246])+$signed(in[157])+$signed(in[282])+$signed(in[283])+$signed(in[94])+$signed(in[284])+$signed(in[125])+$signed(in[158])+$signed(-in[408])+$signed(-in[71])+$signed(-in[97])+$signed(-in[49])+$signed(-in[409])+$signed(-in[165])+$signed(-in[50])+$signed(-in[291])+$signed(-in[229])+$signed(-in[485])+$signed(-in[292])+$signed(-in[110])+$signed(-in[149])+$signed(-in[278])+$signed(-in[422])+$signed(-in[279]);
	sharing32_w = $signed({in[64],1'b0})+$signed({in[384],1'b0})+$signed({in[418],1'b0})+$signed({in[387],1'b0})+$signed(in[451])+$signed({in[164],1'b0})+$signed(in[484])+$signed({in[165],1'b0})+$signed({in[389],1'b0})+$signed(in[262])+$signed({in[231],1'b0})+$signed({in[233],1'b0})+$signed(in[73])+$signed(in[74])+$signed(in[235])+$signed({in[397],1'b0})+$signed(in[430])+$signed({in[399],1'b0})+$signed(in[239])+$signed(in[48])+$signed(in[112])+$signed({in[401],1'b0})+$signed(in[370])+$signed({in[51],1'b0})+$signed({in[244],1'b0})+$signed(in[119])+$signed({in[411],1'b0})+$signed(-in[464])+$signed(-in[130])+$signed(-in[354])+$signed(-in[355])+$signed(-{in[188],1'b0})+$signed(-in[476])+$signed(-in[477])+$signed(-in[270])+$signed(-in[85])+$signed(-in[39]);
	sharing33_w = $signed(in[139])+$signed(in[490])+$signed(in[302])+$signed(in[253])+$signed(-in[365])+$signed(-in[66])+$signed(-in[133])+$signed(-in[495])+$signed(-{in[391],1'b0})+$signed(-in[87]);
	sharing34_w = $signed(in[320])+$signed(in[384])+$signed(in[33])+$signed(in[385])+$signed(in[489])+$signed(in[386])+$signed(in[370])+$signed(in[151])+$signed(in[139])+$signed(in[499])+$signed(in[500])+$signed(in[220])+$signed(in[149])+$signed(in[319])+$signed(-in[117])+$signed(-in[416])+$signed(-in[305])+$signed(-in[155])+$signed(-{in[269],1'b0})+$signed(-in[157])+$signed(-{in[270],1'b0});
	sharing35_w = $signed(in[465])+$signed(in[75])+$signed(in[477])+$signed(in[468])+$signed(in[381])+$signed(in[406])+$signed(in[118])+$signed(in[439])+$signed(-in[229])+$signed(-{in[266],1'b0})+$signed(-in[242])+$signed(-in[191]);
	sharing36_w = $signed(in[465])+$signed(in[17])+$signed(in[482])+$signed({in[131],1'b0})+$signed(in[211])+$signed(in[469])+$signed(in[476])+$signed(in[477])+$signed(in[142])+$signed({in[407],1'b0})+$signed(in[239])+$signed(-{in[192],1'b0})+$signed(-{in[233],2'b0})+$signed(-in[353])+$signed(-{in[402],2'b0})+$signed(-in[76])+$signed(-{in[389],2'b0})+$signed(-in[5])+$signed(-{in[70],1'b0})+$signed(-in[77])+$signed(-in[343]);
	sharing37_w = $signed(in[417])+$signed(in[418])+$signed(in[434])+$signed(in[445])+$signed(-in[504])+$signed(-in[65])+$signed(-in[155])+$signed(-in[203])+$signed(-in[252])+$signed(-in[237])+$signed(-in[279]);
	sharing38_w = $signed(in[328])+$signed(in[384])+$signed(in[410])+$signed(in[394])+$signed(in[331])+$signed(in[244])+$signed(in[79])+$signed(-in[72])+$signed(-in[25])+$signed(-in[137])+$signed(-in[223])+$signed(-in[189])+$signed(-in[343]);
	sharing39_w = $signed({in[160],2'b0})+$signed({in[161],2'b0})+$signed({in[162],2'b0})+$signed({in[163],2'b0})+$signed(in[69])+$signed(in[427])+$signed({in[333],1'b0})+$signed({in[496],1'b0})+$signed(in[401])+$signed(in[146])+$signed(in[50])+$signed({in[149],1'b0})+$signed({in[501],1'b0})+$signed({in[151],1'b0})+$signed(in[152])+$signed(in[216])+$signed(in[219])+$signed(in[251])+$signed(in[220])+$signed(-in[472])+$signed(-in[168])+$signed(-in[368])+$signed(-in[465])+$signed(-in[33])+$signed(-in[121])+$signed(-in[473])+$signed(-in[458])+$signed(-in[298])+$signed(-in[466])+$signed(-in[250])+$signed(-in[463])+$signed(-in[285])+$signed(-in[471]);
	sharing40_w = $signed({in[33],1'b0})+$signed(in[409])+$signed(in[33])+$signed(in[58])+$signed(in[394])+$signed({in[395],1'b0})+$signed(in[163])+$signed({in[396],1'b0})+$signed(in[20])+$signed(in[133])+$signed(in[45])+$signed(in[406])+$signed(in[262])+$signed(in[301])+$signed(-in[49])+$signed(-in[218])+$signed(-in[197]);
	sharing41_w = $signed(in[144])+$signed(in[57])+$signed(in[105])+$signed(in[157])+$signed(in[130])+$signed(in[43])+$signed(in[204])+$signed(in[213])+$signed(-in[357])+$signed(-{in[132],1'b0})+$signed(-{in[373],1'b0})+$signed(-in[21])+$signed(-in[479]);
	sharing42_w = $signed(in[32])+$signed(in[405])+$signed({in[466],1'b0})+$signed(in[250])+$signed(in[426])+$signed(in[469])+$signed(in[315])+$signed(in[379])+$signed(in[29])+$signed(in[317])+$signed({in[30],1'b0})+$signed(in[198])+$signed(in[103])+$signed(-in[321])+$signed(-{in[402],2'b0})+$signed(-in[322])+$signed(-in[203])+$signed(-in[77])+$signed(-in[414])+$signed(-{in[415],1'b0});
	sharing43_w = $signed(in[360])+$signed(in[6])+$signed(in[386])+$signed(in[10])+$signed(in[346])+$signed(in[135])+$signed(in[412])+$signed(in[413])+$signed(in[342])+$signed(in[343])+$signed(-{in[80],1'b0})+$signed(-in[377])+$signed(-in[73])+$signed(-in[257])+$signed(-{in[67],1'b0})+$signed(-in[443])+$signed(-{in[244],1'b0})+$signed(-in[292])+$signed(-{in[245],1'b0})+$signed(-in[453])+$signed(-in[262])+$signed(-in[455]);
	sharing44_w = $signed(in[303])+$signed({in[448],1'b0})+$signed(in[288])+$signed({in[441],1'b0})+$signed(in[497])+$signed(in[290])+$signed(in[482])+$signed(in[498])+$signed(in[90])+$signed(in[499])+$signed(in[453])+$signed(in[461])+$signed({in[367],1'b0})+$signed(in[255])+$signed(-in[385])+$signed(-in[57])+$signed(-{in[412],1'b0})+$signed(-in[396])+$signed(-in[77])+$signed(-{in[166],1'b0})+$signed(-in[93]);
	sharing45_w = $signed(in[193])+$signed(in[17])+$signed(in[505])+$signed(in[426])+$signed(in[355])+$signed({in[204],1'b0})+$signed(in[20])+$signed(in[37])+$signed(in[214])+$signed(-in[316])+$signed(-in[305]);
	sharing46_w = $signed({in[464],1'b0})+$signed(in[256])+$signed(in[240])+$signed({in[465],1'b0})+$signed(in[421])+$signed(in[491])+$signed(in[204])+$signed(in[479])+$signed(in[277])+$signed(in[101])+$signed({in[239],1'b0})+$signed(in[95])+$signed(-in[84])+$signed(-in[362])+$signed(-in[15]);
	sharing47_w = $signed(in[202])+$signed(in[155])+$signed(in[123])+$signed(in[167])+$signed(in[444])+$signed(in[159])+$signed(-in[470])+$signed(-in[144])+$signed(-in[359])+$signed(-in[418])+$signed(-in[42])+$signed(-in[442])+$signed(-in[307])+$signed(-in[395])+$signed(-in[125])+$signed(-in[454])+$signed(-in[333])+$signed(-in[295]);
	sharing48_w = $signed(in[392])+$signed(in[240])+$signed({in[121],1'b0})+$signed(in[337])+$signed(in[42])+$signed(in[146])+$signed(in[291])+$signed(in[27])+$signed(in[318])+$signed(in[495])+$signed(-{in[441],1'b0})+$signed(-{in[289],1'b0})+$signed(-in[18])+$signed(-{in[467],1'b0})+$signed(-in[355])+$signed(-in[358])+$signed(-in[199])+$signed(-{in[302],1'b0})+$signed(-in[78])+$signed(-in[479]);
	sharing49_w = $signed(in[466])+$signed({in[257],1'b0})+$signed(-{in[376],1'b0})+$signed(-in[448])+$signed(-in[145])+$signed(-{in[402],1'b0})+$signed(-in[298])+$signed(-in[461])+$signed(-in[252])+$signed(-in[285])+$signed(-in[438]);
	sharing50_w = $signed({in[456],1'b0})+$signed(in[435])+$signed({in[301],1'b0})+$signed(in[45])+$signed({in[118],1'b0})+$signed(in[38])+$signed(in[422])+$signed({in[455],1'b0})+$signed(in[159])+$signed(-{in[264],1'b0})+$signed(-in[192])+$signed(-{in[272],1'b0})+$signed(-in[405])+$signed(-in[393])+$signed(-{in[276],2'b0})+$signed(-in[61])+$signed(-in[142])+$signed(-{in[94],1'b0})+$signed(-in[230]);
	sharing51_w = $signed(in[289])+$signed(in[290])+$signed({in[291],1'b0})+$signed({in[77],1'b0})+$signed(in[166])+$signed(in[447])+$signed(-{in[278],1'b0})+$signed(-in[410])+$signed(-in[424])+$signed(-in[115]);
	sharing52_w = $signed(in[24])+$signed(in[448])+$signed(in[73])+$signed(in[450])+$signed(in[387])+$signed(in[447])+$signed(in[495])+$signed(in[230])+$signed(in[415])+$signed(-{in[17],1'b0})+$signed(-in[194])+$signed(-{in[355],1'b0})+$signed(-in[212])+$signed(-in[228]);
	sharing53_w = $signed({in[64],1'b0})+$signed(in[344])+$signed(in[153])+$signed({in[402],1'b0})+$signed(in[419])+$signed(in[323])+$signed(in[420])+$signed(in[140])+$signed({in[77],1'b0})+$signed(in[413])+$signed(in[310])+$signed(in[215])+$signed(-{in[416],1'b0})+$signed(-{in[65],1'b0})+$signed(-{in[66],1'b0})+$signed(-in[451])+$signed(-in[452])+$signed(-{in[453],1'b0})+$signed(-{in[390],1'b0})+$signed(-in[294])+$signed(-in[103])+$signed(-in[39])+$signed(-in[107])+$signed(-in[429])+$signed(-in[238])+$signed(-in[78])+$signed(-in[463])+$signed(-in[464])+$signed(-in[113])+$signed(-in[377])+$signed(-in[253])+$signed(-in[126]);
	sharing54_w = $signed(in[109])+$signed(in[216])+$signed(in[408])+$signed(in[96])+$signed(in[240])+$signed(in[113])+$signed(in[213])+$signed(in[188])+$signed(in[21])+$signed(in[197])+$signed(in[95])+$signed(-{in[408],2'b0})+$signed(-in[144])+$signed(-{in[145],1'b0})+$signed(-in[482])+$signed(-{in[315],1'b0})+$signed(-{in[428],1'b0})+$signed(-in[44])+$signed(-in[45])+$signed(-in[31]);
	sharing55_w = $signed(in[89])+$signed(in[233])+$signed(in[466])+$signed(in[391])+$signed(in[123])+$signed(in[259])+$signed(in[231])+$signed(-in[16])+$signed(-in[336])+$signed(-in[394])+$signed(-in[155])+$signed(-in[228]);
	sharing56_w = $signed(in[206])+$signed(in[128])+$signed(in[121])+$signed(in[217])+$signed(in[17])+$signed(in[9])+$signed(in[10])+$signed(in[362])+$signed(in[18])+$signed(in[186])+$signed(in[474])+$signed({in[204],1'b0})+$signed({in[188],1'b0})+$signed(in[439])+$signed({in[22],1'b0})+$signed(in[310])+$signed(in[279])+$signed(-in[65])+$signed(-in[503]);
	sharing57_w = $signed({in[144],1'b0})+$signed(in[145])+$signed(in[241])+$signed({in[242],1'b0})+$signed(in[322])+$signed(in[210])+$signed(in[378])+$signed(in[251])+$signed(in[380])+$signed({in[495],1'b0})+$signed(in[255])+$signed(-{in[400],1'b0})+$signed(-{in[415],1'b0})+$signed(-in[290])+$signed(-{in[76],1'b0})+$signed(-in[68])+$signed(-in[388])+$signed(-in[276])+$signed(-in[493])+$signed(-{in[246],1'b0})+$signed(-{in[63],1'b0})+$signed(-in[87]);
	sharing58_w = $signed({in[296],1'b0})+$signed(in[16])+$signed({in[295],1'b0})+$signed({in[458],1'b0})+$signed(in[162])+$signed(in[298])+$signed({in[114],1'b0})+$signed(in[342])+$signed(in[285])+$signed(in[125])+$signed(in[414])+$signed({in[119],1'b0})+$signed(in[383])+$signed(-in[80])+$signed(-in[56])+$signed(-in[98])+$signed(-in[67])+$signed(-in[404])+$signed(-in[277])+$signed(-in[269])+$signed(-in[54])+$signed(-in[69]);
	sharing59_w = $signed(in[48])+$signed({in[290],1'b0})+$signed(in[146])+$signed(in[291])+$signed(in[211])+$signed(in[109])+$signed(in[110])+$signed(in[359])+$signed(-in[240])+$signed(-in[106])+$signed(-in[283])+$signed(-in[100])+$signed(-in[365])+$signed(-in[334])+$signed(-in[271])+$signed(-in[263]);
	sharing60_w = $signed(in[289])+$signed(in[466])+$signed({in[435],1'b0})+$signed(in[451])+$signed(in[203])+$signed(in[189])+$signed(in[447])+$signed(-in[72])+$signed(-in[8])+$signed(-in[365])+$signed(-in[253]);
	sharing61_w = $signed(in[472])+$signed({in[97],2'b0})+$signed({in[449],1'b0})+$signed(in[109])+$signed(in[199])+$signed(-in[39])+$signed(-in[40])+$signed(-in[496])+$signed(-in[248])+$signed(-{in[65],1'b0})+$signed(-in[429])+$signed(-in[59])+$signed(-in[91])+$signed(-in[132])+$signed(-in[52])+$signed(-in[404])+$signed(-in[157])+$signed(-{in[327],1'b0})+$signed(-in[63]);
	sharing62_w = $signed(in[128])+$signed({in[250],1'b0})+$signed(in[82])+$signed({in[410],1'b0})+$signed(in[460])+$signed({in[79],1'b0})+$signed(in[263])+$signed(-in[392])+$signed(-in[496])+$signed(-in[329])+$signed(-in[117])+$signed(-in[22]);
	sharing63_w = $signed({in[420],1'b0})+$signed(in[202])+$signed(in[102])+$signed(in[421])+$signed(-in[336])+$signed(-in[217])+$signed(-in[505])+$signed(-in[106])+$signed(-in[227])+$signed(-in[70])+$signed(-in[493])+$signed(-{in[142],1'b0})+$signed(-in[94])+$signed(-in[47]);
	sharing64_w = $signed(in[335])+$signed({in[505],1'b0})+$signed(in[433])+$signed(in[402])+$signed({in[291],1'b0})+$signed({in[371],1'b0})+$signed(in[245])+$signed(in[28])+$signed(in[60])+$signed(in[492])+$signed(in[165])+$signed(in[230])+$signed(in[93])+$signed(-in[283])+$signed(-in[228])+$signed(-{in[189],1'b0})+$signed(-{in[191],1'b0})+$signed(-in[351]);
	sharing65_w = $signed(in[140])+$signed(in[206])+$signed(in[19])+$signed(-{in[224],1'b0})+$signed(-{in[393],1'b0})+$signed(-in[249])+$signed(-{in[42],1'b0})+$signed(-{in[366],1'b0})+$signed(-in[382]);
	sharing66_w = $signed(in[400])+$signed(in[24])+$signed(in[488])+$signed(in[228])+$signed(in[254])+$signed(-in[304]);
	sharing67_w = $signed(in[97])+$signed(in[289])+$signed(in[34])+$signed(in[371])+$signed(in[267])+$signed(in[62])+$signed(in[134])+$signed(in[438])+$signed(-{in[264],1'b0})+$signed(-in[281])+$signed(-{in[282],1'b0})+$signed(-in[294])+$signed(-{in[283],1'b0})+$signed(-{in[445],1'b0})+$signed(-in[5])+$signed(-in[94]);
	sharing68_w = $signed(in[401])+$signed({in[68],1'b0})+$signed({in[239],1'b0})+$signed(in[69])+$signed(-in[154])+$signed(-in[204]);
	sharing69_w = $signed({in[144],1'b0})+$signed({in[105],1'b0})+$signed({in[481],1'b0})+$signed({in[20],1'b0})+$signed(in[453])+$signed(in[494])+$signed({in[495],1'b0})+$signed(-{in[24],1'b0})+$signed(-{in[417],2'b0})+$signed(-in[189])+$signed(-in[427])+$signed(-in[333])+$signed(-{in[23],1'b0})+$signed(-in[199]);
	sharing70_w = $signed(in[434])+$signed(in[459])+$signed(in[108])+$signed(in[461])+$signed(in[367])+$signed(-in[136])+$signed(-in[400])+$signed(-in[377])+$signed(-in[322])+$signed(-{in[67],1'b0})+$signed(-in[38]);
	sharing71_w = $signed(in[218])+$signed(in[158])+$signed(in[437])+$signed(-in[470])+$signed(-in[32])+$signed(-{in[369],1'b0})+$signed(-in[297])+$signed(-in[18])+$signed(-in[140])+$signed(-in[150])+$signed(-{in[407],1'b0});
	sharing72_w = $signed({in[160],1'b0})+$signed({in[161],1'b0})+$signed(in[393])+$signed(in[92])+$signed({in[93],1'b0})+$signed(in[333])+$signed(in[222])+$signed(in[159])+$signed(-{in[16],1'b0})+$signed(-in[154])+$signed(-in[290])+$signed(-in[505]);
	sharing73_w = $signed(in[71])+$signed(-in[120])+$signed(-{in[211],1'b0})+$signed(-{in[212],1'b0})+$signed(-in[148])+$signed(-in[310])+$signed(-in[103]);
	sharing74_w = $signed(in[200])+$signed(in[440])+$signed(in[56])+$signed({in[89],1'b0})+$signed(in[297])+$signed(in[201])+$signed(in[410])+$signed({in[19],1'b0})+$signed({in[20],1'b0})+$signed({in[380],1'b0})+$signed({in[373],1'b0})+$signed({in[381],1'b0})+$signed(in[294])+$signed({in[31],1'b0})+$signed(in[367])+$signed(-in[431])+$signed(-in[94])+$signed(-in[428])+$signed(-in[243]);
	sharing75_w = $signed(in[145])+$signed(-{in[290],1'b0})+$signed(-in[448])+$signed(-in[139]);
	sharing76_w = $signed({in[200],1'b0})+$signed(in[192])+$signed(in[280])+$signed(in[153])+$signed(in[217])+$signed(in[130])+$signed(in[122])+$signed(in[322])+$signed(in[187])+$signed(in[476])+$signed(in[486])+$signed(in[463])+$signed(-{in[164],1'b0})+$signed(-in[389])+$signed(-{in[423],1'b0})+$signed(-in[495]);
	sharing77_w = $signed(in[320])+$signed(in[432])+$signed(in[151])+$signed(in[150])+$signed(in[31])+$signed(-in[272])+$signed(-in[81])+$signed(-in[5])+$signed(-{in[430],1'b0})+$signed(-in[46])+$signed(-{in[79],1'b0});
	sharing78_w = $signed(in[464])+$signed(in[56])+$signed(in[129])+$signed(in[107])+$signed(in[380])+$signed(in[382])+$signed(in[302])+$signed(-{in[427],1'b0})+$signed(-in[423]);
	sharing79_w = $signed(in[344])+$signed(in[233])+$signed(in[377])+$signed(in[402])+$signed(in[20])+$signed(in[236])+$signed(in[93])+$signed(in[471])+$signed(-in[420])+$signed(-in[265])+$signed(-in[23]);
	sharing80_w = $signed({in[402],1'b0})+$signed({in[51],1'b0})+$signed(in[123])+$signed({in[220],1'b0})+$signed(in[141])+$signed({in[374],1'b0})+$signed(in[190])+$signed({in[375],1'b0})+$signed(-in[369])+$signed(-in[379])+$signed(-in[403])+$signed(-in[78])+$signed(-in[79]);
	sharing81_w = $signed(in[74])+$signed(in[356])+$signed(in[83])+$signed(in[359])+$signed(-in[280])+$signed(-in[480])+$signed(-in[441])+$signed(-in[482])+$signed(-in[142]);
	sharing82_w = $signed(in[101])+$signed({in[496],1'b0})+$signed({in[160],1'b0})+$signed(in[104])+$signed({in[328],1'b0})+$signed(in[377])+$signed(in[250])+$signed(in[197])+$signed(in[237])+$signed(in[236])+$signed(in[389])+$signed({in[446],1'b0})+$signed({in[167],1'b0})+$signed(in[119])+$signed(-in[480])+$signed(-{in[106],2'b0})+$signed(-in[154])+$signed(-in[491])+$signed(-in[373]);
	sharing83_w = $signed(in[453])+$signed(in[71])+$signed(-in[324]);
	sharing84_w = $signed(in[72])+$signed(in[304])+$signed(in[449])+$signed(in[302])+$signed(in[219])+$signed(in[84])+$signed(in[436])+$signed(in[254])+$signed(-in[363])+$signed(-in[351]);
	sharing85_w = $signed(in[56])+$signed(in[424])+$signed(in[425])+$signed(in[402])+$signed(in[250])+$signed({in[389],1'b0})+$signed(in[437])+$signed(in[446])+$signed(-in[105])+$signed(-in[289])+$signed(-in[210])+$signed(-{in[211],1'b0})+$signed(-in[243]);
	sharing86_w = $signed(in[464])+$signed(in[278])+$signed(-{in[142],1'b0})+$signed(-in[422])+$signed(-{in[77],1'b0})+$signed(-in[303]);
	sharing87_w = $signed(in[232])+$signed({in[201],1'b0})+$signed(in[17])+$signed(in[34])+$signed({in[203],1'b0})+$signed(in[51])+$signed({in[212],1'b0})+$signed({in[205],1'b0})+$signed({in[453],1'b0})+$signed(in[190])+$signed({in[103],1'b0})+$signed(in[375])+$signed(-{in[386],1'b0})+$signed(-in[415])+$signed(-{in[385],1'b0})+$signed(-in[159]);
	sharing88_w = $signed(in[309])+$signed(in[488])+$signed(in[321])+$signed(in[127])+$signed(-in[232])+$signed(-in[100])+$signed(-{in[77],1'b0});
	sharing89_w = $signed({in[16],1'b0})+$signed({in[72],1'b0})+$signed(in[353])+$signed(in[393])+$signed(in[436])+$signed({in[189],1'b0})+$signed(in[5])+$signed(in[374])+$signed(in[366])+$signed(in[422])+$signed(-in[357])+$signed(-{in[467],1'b0})+$signed(-in[323])+$signed(-in[397])+$signed(-in[383]);
	sharing90_w = $signed(in[217])+$signed(in[321])+$signed(in[50])+$signed({in[36],1'b0})+$signed({in[140],1'b0})+$signed(in[308])+$signed({in[484],1'b0})+$signed({in[309],1'b0})+$signed({in[22],1'b0})+$signed(in[494])+$signed({in[486],1'b0})+$signed(in[31])+$signed(-in[288])+$signed(-in[257])+$signed(-{in[65],1'b0})+$signed(-in[255]);
	sharing91_w = $signed({in[202],1'b0})+$signed(in[475])+$signed(in[355])+$signed(in[476])+$signed({in[493],1'b0})+$signed(in[302])+$signed({in[303],1'b0});
	sharing92_w = $signed(in[164])+$signed(in[407])+$signed(-in[115])+$signed(-in[101])+$signed(-in[309])+$signed(-in[118])+$signed(-in[127]);
	sharing93_w = $signed({in[480],1'b0})+$signed(in[8])+$signed(in[191])+$signed(in[5])+$signed(in[7])+$signed(-in[289])+$signed(-in[42])+$signed(-in[491])+$signed(-in[275])+$signed(-in[500])+$signed(-in[29])+$signed(-in[231]);
	sharing94_w = $signed({in[105],1'b0})+$signed(in[281])+$signed(in[401])+$signed(in[458])+$signed(in[211])+$signed(in[99])+$signed(in[92])+$signed({in[470],1'b0})+$signed(in[382])+$signed({in[119],1'b0})+$signed(-{in[426],1'b0})+$signed(-{in[427],2'b0})+$signed(-in[267]);
	sharing95_w = $signed(in[235])+$signed(in[102])+$signed({in[75],1'b0})+$signed(in[293])+$signed(-in[134])+$signed(-in[135]);
	sharing96_w = $signed({in[152],1'b0})+$signed({in[385],2'b0})+$signed({in[386],1'b0})+$signed({in[372],1'b0})+$signed(in[423])+$signed(-in[10])+$signed(-in[6]);
	sharing97_w = $signed(in[412])+$signed(in[422])+$signed({in[77],1'b0})+$signed(in[493])+$signed(-in[258])+$signed(-in[468])+$signed(-in[86])+$signed(-in[369]);
	sharing98_w = $signed({in[392],1'b0})+$signed(in[328])+$signed(in[232])+$signed({in[393],1'b0})+$signed(-in[207])+$signed(-in[335]);
	sharing99_w = $signed({in[18],1'b0})+$signed({in[369],1'b0})+$signed(in[355])+$signed(-{in[240],1'b0})+$signed(-in[58]);
	sharing100_w = $signed(in[209])+$signed(in[378])+$signed(in[162])+$signed(in[106])+$signed(in[498])+$signed(in[219])+$signed(in[499])+$signed({in[38],1'b0})+$signed(-in[272])+$signed(-in[90])+$signed(-in[465]);
	sharing101_w = $signed(in[471])+$signed(in[201])+$signed(-in[128]);
	sharing102_w = $signed(in[329])+$signed(in[277])+$signed(in[145]);
	sharing103_w = $signed(in[431])+$signed(in[416])+$signed({in[165],2'b0})+$signed(in[51]);
	sharing104_w = $signed({in[32],1'b0})+$signed(in[65])+$signed(in[114])+$signed(in[398])+$signed(in[430])+$signed({in[31],1'b0})+$signed(-in[361])+$signed(-in[141]);
	sharing105_w = $signed(in[496])+$signed(in[458])+$signed(in[250])+$signed(in[444])+$signed(in[284])+$signed(-in[140])+$signed(-in[224])+$signed(-in[137]);
	sharing106_w = $signed(in[366])+$signed(in[385])+$signed(in[496])+$signed(in[265]);
	sharing107_w = $signed(in[416])+$signed(in[486])+$signed({in[409],1'b0})+$signed(in[298])+$signed({in[395],1'b0})+$signed({in[133],1'b0})+$signed(in[390])+$signed(-in[504])+$signed(-in[226])+$signed(-in[83])+$signed(-in[460])+$signed(-in[246])+$signed(-in[207]);
	sharing108_w = $signed(in[464])+$signed(in[97])+$signed(in[30])+$signed(in[420])+$signed(in[406])+$signed(in[142])+$signed(-in[284])+$signed(-in[455]);
	sharing109_w = $signed(in[365])+$signed(in[225])+$signed({in[267],1'b0})+$signed(in[213])+$signed(in[335])+$signed(-in[161])+$signed(-in[120])+$signed(-in[162])+$signed(-in[417]);
	sharing110_w = $signed({in[480],1'b0})+$signed({in[466],1'b0})+$signed(in[506])+$signed(in[139])+$signed(in[276])+$signed({in[93],1'b0})+$signed(in[238])+$signed(in[311])+$signed(-{in[425],1'b0})+$signed(-in[75])+$signed(-{in[84],1'b0})+$signed(-{in[413],1'b0})+$signed(-in[295]);
	sharing111_w = $signed(in[198])+$signed(in[224])+$signed(-in[444]);
	sharing112_w = $signed(in[456])+$signed({in[35],1'b0})+$signed({in[20],1'b0})+$signed(in[44])+$signed(in[116])+$signed({in[21],1'b0})+$signed(-in[429])+$signed(-{in[66],1'b0})+$signed(-in[91])+$signed(-{in[53],1'b0})+$signed(-in[445]);
	sharing113_w = $signed(in[431])+$signed(-in[311])+$signed(-{in[315],1'b0})+$signed(-in[71]);
	sharing114_w = $signed(in[144])+$signed(in[460])+$signed({in[469],1'b0})+$signed(in[365])+$signed({in[158],1'b0})+$signed({in[495],1'b0})+$signed(-in[503])+$signed(-in[473])+$signed(-in[199]);
	sharing115_w = $signed(in[83])+$signed(in[309])+$signed(-in[265])+$signed(-in[506])+$signed(-{in[275],1'b0})+$signed(-{in[403],1'b0})+$signed(-in[231]);
	sharing116_w = $signed({in[432],1'b0})+$signed({in[434],1'b0})+$signed(in[280])+$signed(in[423])+$signed(-in[25]);
	sharing117_w = $signed(in[160])+$signed(in[428])+$signed(-in[116])+$signed(-in[259])+$signed(-in[118])+$signed(-in[367]);
	sharing118_w = $signed(in[305])+$signed(in[441])+$signed(in[465])+$signed(in[289])+$signed(in[290])+$signed(in[467])+$signed(in[365])+$signed(in[293])+$signed(in[263])+$signed(-in[310]);
	sharing119_w = $signed(in[124])+$signed(in[215])+$signed(-{in[164],1'b0})+$signed(-in[480])+$signed(-{in[495],1'b0})+$signed(-{in[158],1'b0});
	sharing120_w = $signed(in[462])+$signed(in[426])+$signed({in[253],1'b0})+$signed(in[245])+$signed(in[110])+$signed(in[438])+$signed(-in[43])+$signed(-in[396])+$signed(-in[7]);
	sharing121_w = $signed({in[456],1'b0})+$signed(in[497])+$signed({in[482],1'b0})+$signed(in[442])+$signed({in[469],1'b0})+$signed(in[53])+$signed(in[6])+$signed(in[15])+$signed(-{in[233],1'b0});
	sharing122_w = $signed(in[22])+$signed(in[402])+$signed(in[318])+$signed(-{in[256],1'b0})+$signed(-in[440])+$signed(-in[66])+$signed(-{in[268],1'b0})+$signed(-in[86])+$signed(-in[87]);
	sharing123_w = $signed(in[82])+$signed(in[474])+$signed({in[293],1'b0})+$signed(in[124])+$signed(-in[278])+$signed(-in[232]);
	sharing124_w = $signed({in[292],1'b0})+$signed(in[478])+$signed(in[242])+$signed(in[303])+$signed(-in[115])+$signed(-in[222])+$signed(-in[246])+$signed(-in[501]);
	sharing125_w = $signed({in[461],1'b0})+$signed(in[376])+$signed({in[447],1'b0})+$signed(-in[313])+$signed(-in[330])+$signed(-in[331]);
	sharing126_w = $signed(in[396])+$signed({in[166],1'b0})+$signed(in[158])+$signed(in[267])+$signed(-in[168])+$signed(-{in[217],1'b0})+$signed(-{in[219],2'b0})+$signed(-{in[220],2'b0})+$signed(-{in[206],1'b0})+$signed(-{in[415],2'b0})+$signed(-{in[439],1'b0});
	sharing127_w = $signed(in[192])+$signed(in[408])+$signed(in[388])+$signed(in[497])+$signed(-{in[368],1'b0})+$signed(-{in[394],1'b0})+$signed(-in[357]);
	sharing128_w = $signed(in[49])+$signed(in[248])+$signed(in[265])+$signed(in[367])+$signed(-in[395]);
	sharing129_w = $signed(in[426])+$signed(in[331])+$signed(in[43])+$signed(in[396])+$signed(in[36])+$signed(-in[200])+$signed(-in[112])+$signed(-in[459]);
	sharing130_w = $signed(in[290])+$signed({in[467],1'b0})+$signed(in[245])+$signed(-in[410])+$signed(-in[422])+$signed(-in[316]);
	sharing131_w = $signed({in[41],1'b0})+$signed(in[329])+$signed({in[75],1'b0})+$signed({in[163],1'b0})+$signed(in[331])+$signed(in[236])+$signed({in[213],1'b0});
	sharing132_w = $signed(in[503])+$signed(in[398])+$signed(in[296])+$signed(in[227]);
	sharing133_w = $signed(in[92])+$signed(in[157])+$signed(-{in[476],1'b0})+$signed(-in[436])+$signed(-{in[475],1'b0})+$signed(-{in[453],1'b0});
	sharing134_w = $signed({in[482],1'b0})+$signed(in[137])+$signed(in[483])+$signed(-in[256])+$signed(-in[75]);
	sharing135_w = $signed({in[472],1'b0})+$signed(in[136])+$signed({in[259],1'b0})+$signed({in[21],1'b0})+$signed(in[470])+$signed(in[359])+$signed(-{in[64],1'b0});
	sharing136_w = $signed({in[298],1'b0})+$signed({in[490],1'b0})+$signed({in[491],1'b0})+$signed({in[140],1'b0})+$signed({in[477],1'b0})+$signed({in[502],1'b0})+$signed(in[279])+$signed(-in[104]);
	sharing137_w = $signed({in[450],1'b0})+$signed(in[98])+$signed(-in[443])+$signed(-{in[167],1'b0})+$signed(-in[239]);
	sharing138_w = $signed(in[39])+$signed(in[16])+$signed({in[441],1'b0})+$signed(in[156])+$signed(in[468])+$signed(in[103])+$signed(-in[342])+$signed(-in[334])+$signed(-in[424])+$signed(-in[187]);
	sharing139_w = $signed(in[412])+$signed(in[244])+$signed(in[387])+$signed(-in[131])+$signed(-in[151]);
	sharing140_w = $signed(in[88])+$signed({in[36],1'b0})+$signed(in[454])+$signed(-{in[327],1'b0})+$signed(-in[377]);
	sharing141_w = $signed({in[402],1'b0})+$signed(in[457])+$signed(-{in[416],1'b0})+$signed(-in[270])+$signed(-in[380]);
	sharing142_w = $signed(-{in[121],2'b0})+$signed(-{in[465],1'b0})+$signed(-in[218])+$signed(-in[323])+$signed(-in[123])+$signed(-{in[492],1'b0})+$signed(-in[303]);
	sharing143_w = $signed({in[275],1'b0})+$signed({in[265],1'b0})+$signed(in[351])+$signed(-in[381]);
	sharing144_w = $signed(in[392])+$signed(in[449])+$signed(in[446])+$signed(in[373])+$signed(-{in[311],1'b0})+$signed(-in[499]);
	sharing145_w = $signed({in[23],1'b0})+$signed(in[35])+$signed(-in[105]);
	sharing146_w = $signed(in[41])+$signed(in[146])+$signed({in[147],1'b0})+$signed({in[148],1'b0})+$signed({in[485],1'b0})+$signed(in[135])+$signed(-in[100])+$signed(-in[111]);
	sharing147_w = $signed(in[258])+$signed(in[28])+$signed(in[302])+$signed(in[21])+$signed(-{in[258],2'b0})+$signed(-in[69]);
	sharing148_w = $signed(in[463])+$signed(in[193])+$signed(-in[386])+$signed(-in[282]);
	sharing149_w = $signed(in[464])+$signed({in[241],1'b0})+$signed({in[362],1'b0})+$signed(in[266])+$signed({in[71],1'b0})+$signed(in[343])+$signed(-in[230]);
	sharing150_w = $signed(in[246])+$signed(in[37])+$signed(-in[344])+$signed(-in[90])+$signed(-in[315]);
	sharing151_w = $signed({in[58],1'b0})+$signed(in[268])+$signed({in[228],1'b0})+$signed(-in[390])+$signed(-in[34]);
	sharing152_w = $signed({in[376],1'b0})+$signed(in[68])+$signed(in[411])+$signed(-in[470]);
	sharing153_w = $signed(in[146])+$signed(in[106])+$signed(in[114])+$signed(in[62]);
	sharing154_w = $signed({in[446],1'b0})+$signed(in[87])+$signed({in[443],1'b0})+$signed(in[269])+$signed(-in[487]);
	sharing155_w = $signed({in[220],1'b0})+$signed({in[419],1'b0})+$signed(in[81])+$signed(-{in[378],1'b0})+$signed(-in[496]);
	sharing156_w = $signed({in[94],1'b0})+$signed({in[251],1'b0})+$signed(-in[64])+$signed(-in[65])+$signed(-{in[427],1'b0})+$signed(-in[242]);
	sharing157_w = $signed(in[186])+$signed(in[433])+$signed(-in[151]);
	sharing158_w = $signed({in[158],2'b0})+$signed(in[386])+$signed({in[159],1'b0})+$signed(in[397])+$signed(-in[152])+$signed(-{in[489],1'b0})+$signed(-{in[223],1'b0})+$signed(-{in[214],1'b0})+$signed(-{in[215],1'b0});
	sharing159_w = $signed(in[121])+$signed({in[188],1'b0})+$signed(in[354])+$signed(in[363])+$signed(-{in[422],1'b0})+$signed(-in[38])+$signed(-{in[233],1'b0});
	sharing160_w = $signed({in[408],1'b0})+$signed(in[424])+$signed(-{in[92],1'b0});
	sharing161_w = $signed(in[432])+$signed(in[288])+$signed(in[447])+$signed(in[389])+$signed(in[159])+$signed(-in[24]);
	sharing162_w = $signed(in[472])+$signed(-{in[246],1'b0})+$signed(-{in[263],1'b0});
	sharing163_w = $signed(-in[371])+$signed(-in[216])+$signed(-in[157])+$signed(-in[113]);
	sharing164_w = $signed({in[49],1'b0})+$signed({in[425],1'b0})+$signed({in[426],1'b0})+$signed({in[218],1'b0})+$signed({in[412],1'b0})+$signed(in[372])+$signed({in[37],1'b0})+$signed({in[62],1'b0})+$signed(-in[102])+$signed(-in[277]);
	sharing165_w = $signed(in[72])+$signed(in[190])+$signed({in[93],1'b0})+$signed(in[327])+$signed(-{in[298],1'b0})+$signed(-{in[285],1'b0})+$signed(-in[153]);
	sharing166_w = $signed(in[202])+$signed(in[226])+$signed(-{in[288],1'b0})+$signed(-in[378])+$signed(-in[117]);
	sharing167_w = $signed(in[481])+$signed(-{in[284],1'b0})+$signed(-in[52])+$signed(-in[307])+$signed(-in[101]);
	sharing168_w = $signed({in[50],1'b0})+$signed(in[27])+$signed(-{in[384],1'b0})+$signed(-in[330])+$signed(-in[420])+$signed(-{in[397],1'b0})+$signed(-{in[383],2'b0});
	sharing169_w = $signed(in[412])+$signed(in[168])+$signed(in[501])+$signed(-in[264])+$signed(-in[404])+$signed(-in[130]);
	sharing170_w = $signed(in[489])+$signed(in[283])+$signed({in[103],1'b0})+$signed(in[263]);
	sharing171_w = $signed(in[437])+$signed(in[21])+$signed(-in[66]);
	sharing172_w = $signed(in[154])+$signed(in[424])+$signed({in[203],1'b0})+$signed(in[201])+$signed(-{in[88],1'b0})+$signed(-in[420])+$signed(-in[81]);
	sharing173_w = $signed(in[268])+$signed(in[204])+$signed(in[288])+$signed(in[124])+$signed(-in[117]);
	sharing174_w = $signed({in[402],1'b0})+$signed(in[449])+$signed(in[291]);
	sharing175_w = $signed({in[418],2'b0})+$signed(in[235])+$signed(-in[96])+$signed(-in[457]);
	sharing176_w = $signed({in[242],1'b0})+$signed(-{in[22],1'b0})+$signed(-{in[401],1'b0})+$signed(-in[21]);
	sharing177_w = $signed(in[386])+$signed(-in[43])+$signed(-in[138])+$signed(-{in[379],1'b0})+$signed(-in[53]);
	sharing178_w = $signed({in[456],1'b0})+$signed({in[131],1'b0})+$signed(-in[142]);
	sharing179_w = $signed(in[491])+$signed(in[150])+$signed(in[163])+$signed(-in[252]);
	sharing180_w = $signed({in[370],1'b0})+$signed({in[236],1'b0})+$signed({in[396],1'b0})+$signed(-in[10])+$signed(-in[227]);
	sharing181_w = $signed(in[266])+$signed(in[376])+$signed(in[257]);
	sharing182_w = $signed({in[434],1'b0})+$signed(in[29])+$signed({in[437],1'b0})+$signed(in[101])+$signed(in[407])+$signed(-{in[504],1'b0})+$signed(-in[337]);
	sharing183_w = $signed(in[384])+$signed(in[292])+$signed(in[461])+$signed(-{in[18],2'b0})+$signed(-{in[199],1'b0});
	sharing184_w = $signed({in[430],1'b0})+$signed(in[248])+$signed(in[79])+$signed(-in[321]);
	sharing185_w = $signed(in[160])+$signed(in[345])+$signed(-in[311]);
	sharing186_w = $signed(in[241])+$signed(in[475])+$signed(-in[74])+$signed(-{in[335],1'b0})+$signed(-in[153]);
	sharing187_w = $signed({in[440],1'b0})+$signed(in[53])+$signed(-in[47]);
	sharing188_w = $signed({in[468],1'b0})+$signed(in[332])+$signed({in[479],1'b0})+$signed(in[506]);
	sharing189_w = $signed(in[80])+$signed(in[304])+$signed(-in[28])+$signed(-{in[433],2'b0});
	sharing190_w = $signed({in[189],1'b0})+$signed(-in[71])+$signed(-in[55]);
	sharing191_w = $signed({in[354],1'b0})+$signed(in[202])+$signed({in[357],1'b0})+$signed(in[122])+$signed(-{in[158],1'b0});
	sharing192_w = $signed(in[77])+$signed(-{in[280],1'b0})+$signed(-in[187])+$signed(-{in[281],1'b0})+$signed(-in[39]);
	sharing193_w = $signed(in[126])+$signed({in[375],1'b0})+$signed(-in[72])+$signed(-{in[417],1'b0})+$signed(-in[105]);
	sharing194_w = $signed(in[97])+$signed(in[228])+$signed(in[215])+$signed(in[427])+$signed(-in[164])+$signed(-in[67]);
	sharing195_w = $signed(-in[262])+$signed(-in[226])+$signed(-in[93]);
	sharing196_w = $signed(in[205])+$signed({in[471],1'b0})+$signed(in[133]);
	sharing197_w = $signed({in[461],1'b0})+$signed(-in[436])+$signed(-in[89]);
	sharing198_w = $signed(in[346])+$signed(in[336])+$signed(in[64])+$signed(in[433])+$signed(-in[61]);
	sharing199_w = $signed(in[125])+$signed(-in[212])+$signed(-in[48])+$signed(-in[375]);
	sharing200_w = $signed(in[237])+$signed(in[425])+$signed(-in[119]);
	sharing201_w = $signed(in[240])+$signed({in[154],1'b0})+$signed({in[323],1'b0})+$signed({in[324],1'b0})+$signed({in[141],1'b0})+$signed(-in[76])+$signed(-in[363]);
	sharing202_w = $signed({in[259],1'b0})+$signed({in[359],1'b0})+$signed(in[25])+$signed(-in[199]);
	sharing203_w = $signed(in[223])+$signed(-in[289])+$signed(-in[271])+$signed(-in[115]);
	sharing204_w = $signed(in[78])+$signed(in[77])+$signed({in[495],1'b0})+$signed(in[63])+$signed(-{in[20],2'b0})+$signed(-in[188]);
	sharing205_w = $signed(in[8])+$signed(-in[110])+$signed(-{in[503],1'b0});
	sharing206_w = $signed({in[238],1'b0})+$signed(in[60])+$signed(in[193])+$signed(in[318])+$signed(-{in[64],1'b0})+$signed(-in[356]);
	sharing207_w = $signed(in[164])+$signed(-in[445])+$signed(-in[91]);
	sharing208_w = $signed(in[9])+$signed(-{in[114],1'b0})+$signed(-in[450]);
	sharing209_w = $signed(in[132])+$signed(in[492])+$signed({in[389],1'b0})+$signed(-in[254]);
	sharing210_w = $signed(in[131])+$signed(in[485])+$signed(-{in[458],1'b0})+$signed(-in[212])+$signed(-in[358])+$signed(-in[372]);
	sharing211_w = $signed(in[276])+$signed(in[403])+$signed(-in[295])+$signed(-in[285]);
	sharing212_w = $signed({in[303],1'b0})+$signed({in[159],1'b0})+$signed(-in[418]);
	sharing213_w = $signed(in[86])+$signed(-in[80])+$signed(-in[263]);
	sharing214_w = $signed({in[250],1'b0})+$signed(in[306])+$signed(in[249])+$signed(-in[478]);
	sharing215_w = $signed(in[389])+$signed(-{in[74],1'b0})+$signed(-in[370])+$signed(-in[313]);
	sharing216_w = $signed(in[452])+$signed(-in[287])+$signed(-in[89]);
	sharing217_w = $signed({in[336],1'b0})+$signed(in[502])+$signed({in[289],1'b0})+$signed({in[63],1'b0})+$signed(-in[212])+$signed(-in[116]);
	sharing218_w = $signed({in[230],1'b0})+$signed({in[497],1'b0})+$signed(in[147])+$signed(-{in[454],2'b0})+$signed(-{in[129],2'b0})+$signed(-{in[103],2'b0});
	sharing219_w = $signed({in[417],1'b0})+$signed(-{in[488],1'b0})+$signed(-{in[372],1'b0})+$signed(-{in[487],1'b0});
	sharing220_w = $signed({in[202],1'b0})+$signed(in[465])+$signed(in[319])+$signed(-{in[470],1'b0});
	sharing221_w = $signed(in[459])+$signed(in[391])+$signed(-{in[391],2'b0});
	sharing222_w = $signed({in[50],2'b0})+$signed(in[444])+$signed(in[253]);
	sharing223_w = $signed(in[454])+$signed(in[37])+$signed(-{in[454],2'b0})+$signed(-{in[263],2'b0});
	sharing224_w = $signed({in[114],1'b0})+$signed(-in[18])+$signed(-in[438]);
	sharing225_w = $signed(in[204])+$signed(in[283])+$signed(in[81])+$signed(-in[163]);
	sharing226_w = $signed({in[118],1'b0})+$signed(in[327])+$signed(-{in[64],2'b0});
	sharing227_w = $signed(in[32])+$signed(in[504])+$signed(-in[225]);
	sharing228_w = $signed(in[272])+$signed(in[332])+$signed(in[251])+$signed(-in[132])+$signed(-in[73]);
	sharing229_w = $signed(in[469])+$signed({in[493],1'b0})+$signed(in[59])+$signed(-{in[365],1'b0});
	sharing230_w = $signed(in[36])+$signed(-in[306])+$signed(-in[413]);
	sharing231_w = $signed(in[294])+$signed(in[428])+$signed(in[308])+$signed(-in[25]);
	sharing232_w = $signed({in[66],1'b0})+$signed({in[249],1'b0})+$signed(-in[493]);
	sharing233_w = $signed(-{in[264],1'b0})+$signed(-{in[272],1'b0})+$signed(-{in[465],1'b0})+$signed(-{in[403],2'b0})+$signed(-{in[276],2'b0});
	sharing234_w = $signed({in[216],1'b0})+$signed(in[236])+$signed(in[19])+$signed(-{in[398],1'b0})+$signed(-{in[399],1'b0});
	sharing235_w = $signed(in[102])+$signed(in[191])+$signed(-{in[454],1'b0})+$signed(-in[373]);
	sharing236_w = $signed({in[410],1'b0})+$signed({in[443],1'b0})+$signed(in[487]);
	sharing237_w = $signed(in[466])+$signed({in[371],1'b0})+$signed(in[359]);
	sharing238_w = $signed(in[421])+$signed(in[320])+$signed(in[95])+$signed(-{in[236],1'b0});
	sharing239_w = $signed(in[214])+$signed(-in[333])+$signed(-in[61]);
	sharing240_w = $signed(in[401])+$signed(in[297])+$signed(-in[92]);
	sharing241_w = $signed({in[398],2'b0})+$signed(-{in[200],1'b0})+$signed(-in[210]);
	sharing242_w = $signed(in[485])+$signed(in[410])+$signed(in[220])+$signed(in[55]);
	sharing243_w = $signed(-{in[30],2'b0})+$signed(-in[482])+$signed(-{in[202],2'b0});
	sharing244_w = $signed(in[385])+$signed({in[427],1'b0})+$signed(in[233]);
	sharing245_w = $signed(in[381])+$signed({in[301],1'b0})+$signed(in[111]);
	sharing246_w = $signed({in[322],1'b0})+$signed(in[138])+$signed({in[153],1'b0})+$signed(-in[379]);
	sharing247_w = $signed({in[110],2'b0})+$signed({in[460],1'b0})+$signed(in[467])+$signed(-{in[378],1'b0});
	sharing248_w = $signed(in[200])+$signed(in[50])+$signed(-in[453]);
	sharing249_w = $signed({in[448],1'b0})+$signed(-in[76])+$signed(-in[65]);
	sharing250_w = $signed({in[83],1'b0})+$signed(-in[309])+$signed(-in[79]);
	sharing251_w = $signed({in[190],1'b0})+$signed({in[192],1'b0})+$signed(in[3])+$signed(-in[430]);
	sharing252_w = $signed({in[139],1'b0})+$signed({in[291],1'b0})+$signed({in[33],1'b0})+$signed(in[127]);
	sharing253_w = $signed(in[411])+$signed(in[187])+$signed(-in[54])+$signed(-in[316]);
	sharing254_w = $signed({in[120],1'b0})+$signed({in[122],1'b0})+$signed(in[161]);
	sharing255_w = $signed(in[362])+$signed(-in[70])+$signed(-in[28]);
end

assign weighted_sum[0] = $signed(-{in[192],2'b0})+$signed(-{in[193],1'b0})+$signed(-in[97])+$signed({in[450],1'b0})+$signed(in[34])+$signed({in[68],1'b0})+$signed({in[420],1'b0})+$signed({in[69],1'b0})+$signed(in[37])+$signed({in[421],1'b0})+$signed(in[359])+$signed({in[232],1'b0})+$signed(-{in[360],1'b0})+$signed(-in[424])+$signed(-{in[361],1'b0})+$signed(-{in[362],1'b0})+$signed(-in[426])+$signed({in[491],1'b0})+$signed(in[141])+$signed(in[142])+$signed(-{in[367],2'b0})+$signed({in[431],1'b0})+$signed(in[303])+$signed({in[432],1'b0})+$signed({in[50],1'b0})+$signed(-{in[20],1'b0})+$signed(-in[52])+$signed(-{in[21],1'b0})+$signed({in[373],1'b0})+$signed({in[405],1'b0})+$signed({in[374],1'b0})+$signed(in[214])+$signed({in[407],1'b0})+$signed(in[151])+$signed(in[375])+$signed(-{in[24],1'b0})+$signed(-in[344])+$signed({in[409],1'b0})+$signed(-in[89])+$signed({in[155],1'b0})+$signed({in[219],1'b0})+$signed(-{in[28],2'b0})+$signed({in[92],1'b0})+$signed(-{in[380],1'b0})+$signed(-{in[29],1'b0})+$signed(-{in[30],1'b0})+$signed(-{in[223],1'b0})+$signed(sharing0_r)+$signed(sharing1_r)+$signed(sharing32_r)+$signed(sharing33_r)+$signed(sharing64_r)+$signed(sharing65_r)+$signed(sharing96_r)+$signed(sharing97_r)+$signed(sharing127_r)+$signed(sharing128_r)+$signed(sharing155_r)+$signed(sharing177_r)+$signed(sharing201_r)+$signed(sharing217_r)+$signed(sharing230_r)+$signed(sharing236_r)+$signed(sharing241_r)+$signed(1);
assign weighted_sum[1] = $signed(in[480])+$signed(-{in[65],2'b0})+$signed({in[129],1'b0})+$signed(in[418])+$signed({in[355],1'b0})+$signed(-{in[100],1'b0})+$signed(-in[452])+$signed(in[484])+$signed(in[486])+$signed(in[6])+$signed(in[38])+$signed(-{in[423],1'b0})+$signed(in[136])+$signed(-in[328])+$signed(-{in[265],1'b0})+$signed({in[138],1'b0})+$signed(in[395])+$signed(-in[268])+$signed(in[45])+$signed(-{in[430],2'b0})+$signed(in[46])+$signed({in[144],1'b0})+$signed({in[308],1'b0})+$signed(in[148])+$signed(-in[53])+$signed(in[309])+$signed(-in[279])+$signed(-in[55])+$signed(in[375])+$signed(-{in[376],1'b0})+$signed(in[408])+$signed({in[89],1'b0})+$signed(-in[253])+$signed(in[126])+$signed(sharing2_r)+$signed(sharing3_r)+$signed(sharing34_r)+$signed(sharing35_r)+$signed(sharing66_r)+$signed(sharing67_r)+$signed(sharing104_r)+$signed(-sharing105_r)+$signed(sharing129_r)+$signed(sharing130_r)+$signed(-sharing165_r)+$signed(sharing178_r)+$signed(sharing179_r)+$signed(sharing202_r)+$signed(-2);
assign weighted_sum[2] = $signed(in[128])+$signed(in[480])+$signed(-{in[418],3'b0})+$signed({in[418],1'b0})+$signed(in[162])+$signed(-{in[67],2'b0})+$signed(-{in[387],1'b0})+$signed(-{in[68],3'b0})+$signed(-{in[388],3'b0})+$signed(-{in[69],3'b0})+$signed(-{in[37],1'b0})+$signed(in[357])+$signed({in[69],1'b0})+$signed(-in[166])+$signed(in[455])+$signed(in[231])+$signed({in[40],1'b0})+$signed(in[104])+$signed({in[41],1'b0})+$signed(-in[361])+$signed({in[394],1'b0})+$signed(in[42])+$signed(-{in[238],2'b0})+$signed(in[46])+$signed(-{in[239],3'b0})+$signed(-{in[79],1'b0})+$signed(-in[175])+$signed({in[367],1'b0})+$signed(-{in[80],2'b0})+$signed(-in[431])+$signed(in[467])+$signed({in[116],1'b0})+$signed(-in[405])+$signed(-{in[406],2'b0})+$signed(-{in[246],1'b0})+$signed(-in[278])+$signed(-{in[407],3'b0})+$signed(-{in[375],2'b0})+$signed(-{in[408],3'b0})+$signed(-{in[56],1'b0})+$signed({in[408],1'b0})+$signed(-{in[57],1'b0})+$signed(-{in[89],1'b0})+$signed({in[442],1'b0})+$signed(-in[186])+$signed(-{in[187],1'b0})+$signed(in[61])+$signed({in[158],1'b0})+$signed(in[94])+$signed(in[127])+$signed(sharing24_r)+$signed(-sharing25_r)+$signed(sharing36_r)+$signed(sharing37_r)+$signed(sharing68_r)+$signed(sharing69_r)+$signed(sharing98_r)+$signed(sharing99_r)+$signed(-sharing155_r)+$signed(sharing180_r)+$signed(sharing226_r)+$signed(-sharing235_r)+$signed(sharing237_r)+$signed(0);
assign weighted_sum[3] = $signed(-in[480])+$signed({in[385],1'b0})+$signed(in[129])+$signed(-in[1])+$signed({in[226],1'b0})+$signed(-in[194])+$signed({in[227],1'b0})+$signed(in[67])+$signed({in[100],1'b0})+$signed(-in[4])+$signed({in[132],1'b0})+$signed({in[388],1'b0})+$signed(in[420])+$signed(-in[358])+$signed({in[424],1'b0})+$signed(-in[168])+$signed(in[457])+$signed(-in[489])+$signed({in[74],1'b0})+$signed(in[234])+$signed(-{in[298],1'b0})+$signed(in[427])+$signed({in[398],1'b0})+$signed(-in[110])+$signed({in[207],1'b0})+$signed(in[431])+$signed({in[80],1'b0})+$signed({in[400],1'b0})+$signed({in[433],1'b0})+$signed(in[145])+$signed({in[146],1'b0})+$signed({in[402],1'b0})+$signed(-{in[466],1'b0})+$signed(-{in[467],2'b0})+$signed(-{in[19],1'b0})+$signed({in[243],1'b0})+$signed(-{in[116],2'b0})+$signed(-in[276])+$signed({in[246],1'b0})+$signed(in[189])+$signed(-in[156])+$signed(-{in[189],2'b0})+$signed(-{in[285],1'b0})+$signed(in[61])+$signed(-in[255])+$signed(sharing4_r)+$signed(sharing5_r)+$signed(sharing32_r)+$signed(-sharing33_r)+$signed(sharing72_r)+$signed(-sharing73_r)+$signed(sharing100_r)+$signed(sharing101_r)+$signed(sharing131_r)+$signed(sharing164_r)+$signed(sharing181_r)+$signed(sharing182_r)+$signed(sharing203_r)+$signed(sharing218_r)+$signed(sharing231_r)+$signed(sharing242_r)+$signed(sharing248_r)+$signed(1);
assign weighted_sum[4] = $signed(-{in[128],2'b0})+$signed(in[385])+$signed({in[159],1'b0})+$signed(-{in[355],1'b0})+$signed({in[164],2'b0})+$signed(in[486])+$signed(-in[134])+$signed(in[391])+$signed(in[232])+$signed(in[488])+$signed(-in[361])+$signed(in[393])+$signed({in[330],1'b0})+$signed(-in[362])+$signed({in[331],1'b0})+$signed({in[332],2'b0})+$signed(-{in[301],1'b0})+$signed(in[45])+$signed(-{in[142],1'b0})+$signed(-in[366])+$signed(-{in[16],2'b0})+$signed(in[144])+$signed({in[498],1'b0})+$signed({in[499],1'b0})+$signed(-{in[116],1'b0})+$signed(in[372])+$signed({in[500],1'b0})+$signed(-{in[21],2'b0})+$signed(-{in[22],2'b0})+$signed({in[150],1'b0})+$signed(in[278])+$signed({in[502],2'b0})+$signed(-{in[119],1'b0})+$signed(in[217])+$signed(in[58])+$signed(-in[378])+$signed(in[379])+$signed(-in[443])+$signed(-{in[477],1'b0})+$signed({in[382],1'b0})+$signed(in[446])+$signed(-{in[479],1'b0})+$signed(sharing0_r)+$signed(-sharing1_r)+$signed(sharing38_r)+$signed(sharing39_r)+$signed(sharing92_r)+$signed(-sharing93_r)+$signed(sharing102_r)+$signed(sharing103_r)+$signed(sharing132_r)+$signed(sharing133_r)+$signed(sharing161_r)+$signed(-sharing191_r)+$signed(sharing204_r)+$signed(sharing218_r)+$signed(sharing238_r)+$signed(1);
assign weighted_sum[5] = $signed({in[192],1'b0})+$signed(-in[481])+$signed(-in[33])+$signed(in[98])+$signed(-{in[483],2'b0})+$signed(-{in[484],1'b0})+$signed(-in[132])+$signed(in[292])+$signed(in[324])+$signed(in[389])+$signed(-in[421])+$signed(in[37])+$signed(-in[72])+$signed(in[328])+$signed(-in[456])+$signed(-{in[393],1'b0})+$signed(-in[488])+$signed(-{in[394],2'b0})+$signed(in[458])+$signed(-in[267])+$signed(-{in[77],2'b0})+$signed({in[239],1'b0})+$signed(-in[368])+$signed(in[82])+$signed(-in[243])+$signed(in[435])+$signed(-{in[149],1'b0})+$signed(-{in[246],2'b0})+$signed(in[86])+$signed(-in[374])+$signed(-{in[55],1'b0})+$signed({in[505],1'b0})+$signed(in[281])+$signed(-in[250])+$signed(-{in[411],2'b0})+$signed(-{in[412],2'b0})+$signed(-{in[381],1'b0})+$signed(in[157])+$signed({in[445],1'b0})+$signed(-{in[382],1'b0})+$signed(-in[254])+$signed(-{in[415],2'b0})+$signed(-{in[223],1'b0})+$signed(sharing4_r)+$signed(-sharing5_r)+$signed(sharing54_r)+$signed(-sharing55_r)+$signed(sharing70_r)+$signed(sharing71_r)+$signed(sharing106_r)+$signed(-sharing107_r)+$signed(sharing145_r)+$signed(-sharing146_r)+$signed(sharing156_r)+$signed(sharing157_r)+$signed(-sharing180_r)+$signed(-sharing232_r)+$signed(-sharing236_r)+$signed(-sharing255_r)+$signed(2);
assign weighted_sum[6] = $signed(-{in[96],2'b0})+$signed({in[416],1'b0})+$signed(-in[448])+$signed(-{in[95],1'b0})+$signed(-in[385])+$signed(in[321])+$signed(-in[98])+$signed(-in[35])+$signed(-in[259])+$signed(in[419])+$signed(-{in[356],1'b0})+$signed(in[68])+$signed(-in[100])+$signed({in[452],1'b0})+$signed(in[390])+$signed(-in[422])+$signed({in[71],1'b0})+$signed(-{in[457],1'b0})+$signed(in[41])+$signed(-{in[266],3'b0})+$signed(-{in[106],2'b0})+$signed({in[266],1'b0})+$signed(-{in[107],2'b0})+$signed(-{in[459],1'b0})+$signed(-{in[108],1'b0})+$signed(-in[461])+$signed(-in[462])+$signed(in[239])+$signed(-{in[435],3'b0})+$signed(-{in[19],1'b0})+$signed(in[275])+$signed(-{in[84],2'b0})+$signed(-in[469])+$signed({in[54],1'b0})+$signed(-{in[278],1'b0})+$signed(-in[310])+$signed(-{in[279],2'b0})+$signed({in[55],1'b0})+$signed(-in[215])+$signed(-in[120])+$signed(in[314])+$signed(-{in[444],1'b0})+$signed(-in[254])+$signed(-{in[447],2'b0})+$signed(-{in[223],1'b0})+$signed(sharing12_r)+$signed(-sharing13_r)+$signed(sharing60_r)+$signed(-sharing61_r)+$signed(sharing78_r)+$signed(-sharing79_r)+$signed(sharing98_r)+$signed(-sharing99_r)+$signed(sharing153_r)+$signed(-sharing154_r)+$signed(sharing170_r)+$signed(-sharing171_r)+$signed(-sharing177_r)+$signed(sharing210_r)+$signed(sharing220_r)+$signed(-sharing248_r)+$signed(2);
assign weighted_sum[7] = $signed(in[96])+$signed(-{in[290],2'b0})+$signed(-{in[258],1'b0})+$signed(in[66])+$signed(-{in[291],2'b0})+$signed(in[260])+$signed(in[292])+$signed(-{in[293],2'b0})+$signed(in[326])+$signed(in[455])+$signed(-{in[457],2'b0})+$signed(-in[105])+$signed(-{in[458],2'b0})+$signed(in[330])+$signed(in[426])+$signed(-{in[459],1'b0})+$signed(-{in[76],1'b0})+$signed(-in[108])+$signed(in[332])+$signed(in[141])+$signed(-in[269])+$signed(in[398])+$signed(-{in[303],3'b0})+$signed({in[431],1'b0})+$signed(-{in[304],3'b0})+$signed({in[304],1'b0})+$signed(in[432])+$signed(-{in[305],2'b0})+$signed(in[307])+$signed(in[500])+$signed(in[149])+$signed(-in[245])+$signed(-in[246])+$signed(in[374])+$signed(-{in[119],2'b0})+$signed(-{in[120],3'b0})+$signed(-{in[121],3'b0})+$signed(-{in[473],2'b0})+$signed(in[249])+$signed(-{in[122],3'b0})+$signed(-{in[474],2'b0})+$signed(in[474])+$signed(-{in[123],2'b0})+$signed({in[315],1'b0})+$signed(in[155])+$signed(in[94])+$signed({in[447],1'b0})+$signed(sharing18_r)+$signed(-sharing19_r)+$signed(sharing48_r)+$signed(-sharing49_r)+$signed(sharing82_r)+$signed(-sharing83_r)+$signed(sharing100_r)+$signed(-sharing101_r)+$signed(sharing134_r)+$signed(-sharing135_r)+$signed(-sharing173_r)+$signed(sharing192_r)+$signed(sharing212_r)+$signed(-sharing213_r)+$signed(sharing254_r)+$signed(2);
assign weighted_sum[8] = $signed(-{in[32],3'b0})+$signed(in[32])+$signed(-{in[33],3'b0})+$signed(in[381])+$signed(-{in[34],2'b0})+$signed({in[162],1'b0})+$signed(-in[322])+$signed(-{in[35],2'b0})+$signed(-{in[483],2'b0})+$signed(-{in[484],2'b0})+$signed(-{in[133],2'b0})+$signed(-{in[485],2'b0})+$signed(-{in[134],1'b0})+$signed(-{in[486],1'b0})+$signed(in[167])+$signed(-{in[200],2'b0})+$signed(in[264])+$signed(-{in[201],2'b0})+$signed(-{in[203],2'b0})+$signed(-in[139])+$signed(-{in[204],2'b0})+$signed(in[44])+$signed(-{in[205],1'b0})+$signed(in[429])+$signed(-{in[366],1'b0})+$signed(-{in[367],2'b0})+$signed({in[79],1'b0})+$signed(-{in[368],2'b0})+$signed(-{in[17],2'b0})+$signed(-{in[369],2'b0})+$signed(in[497])+$signed(-{in[370],2'b0})+$signed(-{in[19],2'b0})+$signed(-{in[371],2'b0})+$signed(in[19])+$signed(in[436])+$signed(-{in[213],2'b0})+$signed(-{in[22],1'b0})+$signed(-in[374])+$signed(-in[503])+$signed(-{in[476],1'b0})+$signed(-{in[29],1'b0})+$signed(in[445])+$signed(in[382])+$signed(-{in[31],3'b0})+$signed({in[383],1'b0})+$signed(in[31])+$signed(sharing6_r)+$signed(sharing7_r)+$signed(sharing40_r)+$signed(sharing41_r)+$signed(sharing72_r)+$signed(sharing73_r)+$signed(sharing104_r)+$signed(sharing105_r)+$signed(sharing139_r)+$signed(-sharing140_r)+$signed(sharing158_r)+$signed(sharing183_r)+$signed(sharing184_r)+$signed(sharing204_r)+$signed(sharing219_r)+$signed(sharing232_r)+$signed(sharing243_r)+$signed(2);
assign weighted_sum[9] = $signed(-in[417])+$signed(in[194])+$signed({in[355],1'b0})+$signed(-in[291])+$signed(in[131])+$signed({in[356],1'b0})+$signed(-in[452])+$signed({in[357],1'b0})+$signed(in[485])+$signed(in[101])+$signed({in[358],1'b0})+$signed({in[134],1'b0})+$signed(-in[104])+$signed(in[425])+$signed({in[394],1'b0})+$signed(in[42])+$signed(-in[106])+$signed(-in[107])+$signed(in[237])+$signed(in[397])+$signed(-in[461])+$signed(in[175])+$signed({in[16],1'b0})+$signed({in[17],1'b0})+$signed(-{in[81],1'b0})+$signed(in[18])+$signed(in[114])+$signed({in[467],1'b0})+$signed(-in[275])+$signed({in[471],1'b0})+$signed(-in[279])+$signed({in[473],1'b0})+$signed(in[25])+$signed(-in[217])+$signed({in[90],1'b0})+$signed(in[282])+$signed({in[474],1'b0})+$signed(-in[219])+$signed({in[285],1'b0})+$signed(sharing8_r)+$signed(sharing9_r)+$signed(sharing42_r)+$signed(sharing43_r)+$signed(sharing74_r)+$signed(sharing75_r)+$signed(sharing106_r)+$signed(sharing107_r)+$signed(sharing134_r)+$signed(sharing135_r)+$signed(sharing159_r)+$signed(sharing160_r)+$signed(sharing185_r)+$signed(sharing186_r)+$signed(sharing205_r)+$signed(-sharing217_r)+$signed(1);
assign weighted_sum[10] = $signed({in[128],1'b0})+$signed(in[480])+$signed({in[129],1'b0})+$signed(in[226])+$signed(in[100])+$signed(-in[132])+$signed(-in[484])+$signed({in[454],1'b0})+$signed(in[487])+$signed(-in[7])+$signed(in[199])+$signed(in[488])+$signed({in[201],1'b0})+$signed(-in[233])+$signed({in[42],1'b0})+$signed({in[203],1'b0})+$signed({in[109],1'b0})+$signed(in[109])+$signed(in[205])+$signed({in[369],1'b0})+$signed(in[114])+$signed({in[467],1'b0})+$signed(in[500])+$signed({in[213],1'b0})+$signed(in[149])+$signed({in[501],1'b0})+$signed({in[23],1'b0})+$signed({in[279],1'b0})+$signed(in[311])+$signed(in[24])+$signed(-in[58])+$signed(in[218])+$signed(in[220])+$signed(in[380])+$signed(in[189])+$signed(in[382])+$signed(sharing10_r)+$signed(sharing11_r)+$signed(sharing44_r)+$signed(sharing45_r)+$signed(sharing76_r)+$signed(sharing77_r)+$signed(sharing108_r)+$signed(sharing109_r)+$signed(sharing136_r)+$signed(sharing137_r)+$signed(-sharing158_r)+$signed(sharing187_r)+$signed(sharing188_r)+$signed(-sharing205_r)+$signed(sharing220_r)+$signed(sharing234_r)+$signed(sharing252_r)+$signed(0);
assign weighted_sum[11] = $signed({in[480],1'b0})+$signed(in[416])+$signed({in[66],1'b0})+$signed({in[259],1'b0})+$signed({in[323],1'b0})+$signed(-{in[419],1'b0})+$signed(in[483])+$signed(-{in[420],1'b0})+$signed(in[4])+$signed(-{in[421],2'b0})+$signed(-in[165])+$signed(in[293])+$signed(-in[326])+$signed(in[134])+$signed({in[263],1'b0})+$signed(-in[168])+$signed(in[329])+$signed(-in[457])+$signed(in[459])+$signed(-{in[428],1'b0})+$signed(in[108])+$signed(-in[396])+$signed({in[492],1'b0})+$signed(-in[77])+$signed(in[206])+$signed(-in[401])+$signed(-{in[402],2'b0})+$signed(-{in[435],2'b0})+$signed(-in[51])+$signed({in[52],1'b0})+$signed(in[244])+$signed(-{in[437],1'b0})+$signed(-{in[118],1'b0})+$signed(-in[54])+$signed(in[278])+$signed({in[190],1'b0})+$signed(-{in[409],1'b0})+$signed(in[154])+$signed({in[93],1'b0})+$signed({in[94],1'b0})+$signed(-{in[415],2'b0})+$signed(sharing12_r)+$signed(sharing13_r)+$signed(sharing46_r)+$signed(sharing47_r)+$signed(sharing76_r)+$signed(-sharing77_r)+$signed(sharing124_r)+$signed(-sharing125_r)+$signed(sharing143_r)+$signed(-sharing144_r)+$signed(sharing159_r)+$signed(-sharing160_r)+$signed(sharing189_r)+$signed(sharing190_r)+$signed(sharing206_r)+$signed(-sharing249_r)+$signed(2);
assign weighted_sum[12] = $signed(-in[63])+$signed(-in[481])+$signed(in[225])+$signed(-{in[388],2'b0})+$signed({in[453],1'b0})+$signed(in[133])+$signed(in[229])+$signed(-{in[422],3'b0})+$signed({in[390],1'b0})+$signed(-{in[455],2'b0})+$signed(-{in[263],2'b0})+$signed(-{in[264],2'b0})+$signed(in[40])+$signed(in[136])+$signed(-in[105])+$signed(-{in[426],1'b0})+$signed(in[267])+$signed(in[12])+$signed(-in[205])+$signed(-{in[430],2'b0})+$signed(in[430])+$signed(-{in[431],3'b0})+$signed(in[303])+$signed(-{in[432],3'b0})+$signed(in[495])+$signed({in[368],1'b0})+$signed(-{in[81],3'b0})+$signed({in[81],1'b0})+$signed(in[369])+$signed(-{in[82],3'b0})+$signed(-{in[401],1'b0})+$signed(in[370])+$signed(-{in[83],3'b0})+$signed(-{in[275],1'b0})+$signed(in[403])+$signed(in[116])+$signed(in[277])+$signed(-in[503])+$signed(-in[88])+$signed(in[410])+$signed(-{in[92],2'b0})+$signed(-{in[93],3'b0})+$signed(-{in[253],2'b0})+$signed(-in[285])+$signed(-{in[94],2'b0})+$signed(in[478])+$signed(-in[190])+$signed(in[383])+$signed(sharing14_r)+$signed(sharing15_r)+$signed(sharing36_r)+$signed(-sharing37_r)+$signed(sharing78_r)+$signed(sharing79_r)+$signed(sharing110_r)+$signed(sharing111_r)+$signed(sharing138_r)+$signed(sharing161_r)+$signed(sharing189_r)+$signed(-sharing190_r)+$signed(sharing216_r)+$signed(-sharing231_r)+$signed(sharing245_r)+$signed(sharing250_r)+$signed(1);
assign weighted_sum[13] = $signed(-{in[65],1'b0})+$signed(-{in[129],1'b0})+$signed(-{in[451],2'b0})+$signed({in[227],1'b0})+$signed(-in[35])+$signed(-in[67])+$signed(-{in[36],2'b0})+$signed(-{in[387],1'b0})+$signed(-in[356])+$signed(-{in[388],2'b0})+$signed(-{in[37],2'b0})+$signed(-{in[452],2'b0})+$signed(-{in[262],1'b0})+$signed(-in[102])+$signed(-in[38])+$signed(in[255])+$signed(-{in[392],2'b0})+$signed(-{in[40],1'b0})+$signed(-{in[41],2'b0})+$signed(-{in[233],2'b0})+$signed(-{in[393],2'b0})+$signed(-{in[42],2'b0})+$signed({in[266],1'b0})+$signed(-{in[427],2'b0})+$signed(-in[235])+$signed(in[46])+$signed(-in[366])+$signed({in[399],1'b0})+$signed(-in[207])+$signed(-{in[464],2'b0})+$signed(-{in[401],2'b0})+$signed(-{in[466],2'b0})+$signed(-{in[211],2'b0})+$signed(-in[115])+$signed(-{in[53],2'b0})+$signed(in[85])+$signed({in[214],1'b0})+$signed(in[503])+$signed(-{in[440],2'b0})+$signed(-in[152])+$signed(in[505])+$signed(-{in[218],1'b0})+$signed(-in[26])+$signed(in[122])+$signed(-in[314])+$signed(-{in[379],2'b0})+$signed({in[506],1'b0})+$signed(-{in[380],3'b0})+$signed(in[380])+$signed(-{in[381],3'b0})+$signed({in[381],1'b0})+$signed(-{in[414],1'b0})+$signed(in[30])+$signed(-{in[63],2'b0})+$signed(in[319])+$signed(sharing16_r)+$signed(sharing17_r)+$signed(sharing48_r)+$signed(sharing49_r)+$signed(sharing86_r)+$signed(-sharing87_r)+$signed(sharing126_r)+$signed(sharing127_r)+$signed(-sharing128_r)+$signed(sharing162_r)+$signed(sharing163_r)+$signed(sharing185_r)+$signed(-sharing186_r)+$signed(sharing207_r)+$signed(sharing208_r)+$signed(sharing221_r)+$signed(-sharing222_r)+$signed(sharing233_r)+$signed(-sharing238_r)+$signed(sharing240_r)+$signed(sharing243_r)+$signed(-1);
assign weighted_sum[14] = $signed(-{in[96],1'b0})+$signed(in[64])+$signed(-in[257])+$signed(in[34])+$signed(-{in[259],2'b0})+$signed(-in[4])+$signed(in[100])+$signed(-in[5])+$signed(in[486])+$signed(-in[390])+$signed(in[167])+$signed(in[40])+$signed(in[232])+$signed(in[328])+$signed(-{in[76],2'b0})+$signed(-{in[108],2'b0})+$signed(-{in[109],3'b0})+$signed({in[109],1'b0})+$signed(-in[429])+$signed(in[368])+$signed(in[496])+$signed({in[433],1'b0})+$signed({in[18],1'b0})+$signed(in[402])+$signed(-{in[277],3'b0})+$signed(-{in[245],1'b0})+$signed({in[277],1'b0})+$signed(-{in[278],3'b0})+$signed(in[29])+$signed(in[22])+$signed(-{in[279],2'b0})+$signed(-in[343])+$signed(-{in[280],2'b0})+$signed(-in[88])+$signed(-{in[89],3'b0})+$signed(in[376])+$signed({in[89],1'b0})+$signed(in[121])+$signed(-{in[90],1'b0})+$signed(-{in[445],2'b0})+$signed(-in[413])+$signed(-{in[446],2'b0})+$signed(-{in[95],2'b0})+$signed(in[223])+$signed(sharing18_r)+$signed(sharing19_r)+$signed(sharing50_r)+$signed(-sharing51_r)+$signed(sharing94_r)+$signed(-sharing95_r)+$signed(sharing116_r)+$signed(-sharing117_r)+$signed(sharing147_r)+$signed(-sharing148_r)+$signed(sharing162_r)+$signed(-sharing163_r)+$signed(sharing196_r)+$signed(-sharing197_r)+$signed(sharing209_r)+$signed(-sharing247_r)+$signed(1);
assign weighted_sum[15] = $signed(in[448])+$signed(-{in[417],2'b0})+$signed(in[34])+$signed(-{in[164],1'b0})+$signed(-in[228])+$signed(-in[388])+$signed({in[421],1'b0})+$signed(-in[229])+$signed(-in[230])+$signed(-in[167])+$signed(-{in[328],2'b0})+$signed(-{in[392],1'b0})+$signed(-{in[488],1'b0})+$signed({in[105],1'b0})+$signed(-{in[329],1'b0})+$signed(-{in[330],2'b0})+$signed(-{in[331],2'b0})+$signed(-in[43])+$signed(in[11])+$signed(-{in[332],1'b0})+$signed(in[462])+$signed(-{in[79],2'b0})+$signed(-{in[80],2'b0})+$signed(-{in[497],2'b0})+$signed(-{in[145],1'b0})+$signed(-in[49])+$signed(in[17])+$signed(-{in[498],2'b0})+$signed(-{in[499],2'b0})+$signed(-in[307])+$signed(-{in[500],2'b0})+$signed(in[52])+$signed(in[245])+$signed(-in[341])+$signed(-{in[150],2'b0})+$signed(-in[502])+$signed(-in[215])+$signed(-in[56])+$signed(-{in[250],2'b0})+$signed({in[90],1'b0})+$signed(-in[442])+$signed(in[124])+$signed(-in[93])+$signed(-{in[159],2'b0})+$signed(-{in[319],1'b0})+$signed(in[415])+$signed(sharing26_r)+$signed(-sharing27_r)+$signed(sharing38_r)+$signed(-sharing39_r)+$signed(sharing70_r)+$signed(-sharing71_r)+$signed(sharing108_r)+$signed(-sharing109_r)+$signed(sharing138_r)+$signed(sharing174_r)+$signed(-sharing175_r)+$signed(sharing199_r)+$signed(-sharing200_r)+$signed(-sharing206_r)+$signed(-sharing225_r)+$signed(0);
assign weighted_sum[16] = $signed({in[64],1'b0})+$signed(-{in[481],1'b0})+$signed(-{in[130],1'b0})+$signed(in[291])+$signed(in[259])+$signed(-in[166])+$signed({in[231],1'b0})+$signed(-in[40])+$signed(in[265])+$signed({in[298],1'b0})+$signed(in[106])+$signed(in[75])+$signed(in[203])+$signed(-in[108])+$signed(in[332])+$signed(in[460])+$signed(-{in[237],1'b0})+$signed(-{in[496],2'b0})+$signed({in[48],1'b0})+$signed(in[16])+$signed(-in[336])+$signed(-in[368])+$signed({in[401],1'b0})+$signed(in[306])+$signed(-{in[404],1'b0})+$signed({in[373],2'b0})+$signed(in[342])+$signed({in[23],1'b0})+$signed(in[471])+$signed({in[473],1'b0})+$signed(-{in[505],1'b0})+$signed({in[219],1'b0})+$signed(-in[60])+$signed({in[413],2'b0})+$signed(in[285])+$signed({in[414],2'b0})+$signed({in[191],1'b0})+$signed(sharing20_r)+$signed(sharing21_r)+$signed(sharing56_r)+$signed(-sharing57_r)+$signed(sharing80_r)+$signed(sharing81_r)+$signed(sharing112_r)+$signed(sharing113_r)+$signed(sharing139_r)+$signed(sharing140_r)+$signed(sharing164_r)+$signed(sharing191_r)+$signed(sharing209_r)+$signed(sharing221_r)+$signed(sharing222_r)+$signed(sharing244_r)+$signed(sharing253_r)+$signed(0);
assign weighted_sum[17] = $signed(-{in[288],1'b0})+$signed(in[224])+$signed(in[222])+$signed(-{in[289],2'b0})+$signed(-in[417])+$signed(-{in[290],3'b0})+$signed({in[290],1'b0})+$signed(-in[354])+$signed(-{in[291],3'b0})+$signed(-in[451])+$signed(-{in[292],3'b0})+$signed({in[292],1'b0})+$signed(-{in[452],1'b0})+$signed(-{in[453],2'b0})+$signed(-{in[262],2'b0})+$signed(-{in[232],1'b0})+$signed(-in[392])+$signed(-{in[107],3'b0})+$signed(-{in[459],3'b0})+$signed(in[459])+$signed(-{in[108],3'b0})+$signed(-{in[460],3'b0})+$signed({in[108],1'b0})+$signed(-{in[109],2'b0})+$signed(in[109])+$signed(-in[493])+$signed(-{in[430],2'b0})+$signed(in[46])+$signed(in[15])+$signed(in[47])+$signed(-in[335])+$signed(in[336])+$signed(-in[464])+$signed(in[210])+$signed(in[434])+$signed(-{in[467],2'b0})+$signed(-{in[277],2'b0})+$signed(in[277])+$signed(-{in[439],1'b0})+$signed(-in[311])+$signed(-{in[440],1'b0})+$signed(-{in[89],2'b0})+$signed(-in[505])+$signed(-{in[122],2'b0})+$signed(-{in[250],2'b0})+$signed(in[442])+$signed(in[91])+$signed(-in[251])+$signed(-in[443])+$signed(-{in[92],1'b0})+$signed(in[316])+$signed(-{in[93],3'b0})+$signed(-{in[444],2'b0})+$signed(-{in[445],1'b0})+$signed(-{in[478],1'b0})+$signed(in[414])+$signed(in[287])+$signed(sharing22_r)+$signed(sharing23_r)+$signed(sharing50_r)+$signed(sharing51_r)+$signed(sharing82_r)+$signed(sharing83_r)+$signed(sharing114_r)+$signed(sharing115_r)+$signed(sharing141_r)+$signed(sharing142_r)+$signed(sharing165_r)+$signed(sharing194_r)+$signed(-sharing195_r)+$signed(sharing210_r)+$signed(sharing223_r)+$signed(sharing224_r)+$signed(sharing249_r)+$signed(0);
assign weighted_sum[18] = $signed(-{in[480],1'b0})+$signed(-in[256])+$signed(in[97])+$signed({in[322],1'b0})+$signed(in[98])+$signed(-{in[102],1'b0})+$signed(-{in[198],1'b0})+$signed(-in[262])+$signed(-in[8])+$signed(-in[296])+$signed(-in[41])+$signed(in[394])+$signed(in[490])+$signed(-{in[235],1'b0})+$signed(in[397])+$signed(-in[270])+$signed(-{in[271],2'b0})+$signed(in[303])+$signed(-in[16])+$signed(in[49])+$signed(-in[177])+$signed(-in[337])+$signed(-{in[466],1'b0})+$signed(-{in[275],2'b0})+$signed(in[435])+$signed({in[85],1'b0})+$signed(in[214])+$signed(in[86])+$signed(in[152])+$signed(in[57])+$signed(-{in[282],1'b0})+$signed(-in[90])+$signed(in[218])+$signed(-{in[283],1'b0})+$signed(in[220])+$signed(-in[125])+$signed(sharing24_r)+$signed(sharing25_r)+$signed(sharing52_r)+$signed(sharing53_r)+$signed(sharing84_r)+$signed(sharing85_r)+$signed(sharing116_r)+$signed(sharing117_r)+$signed(sharing129_r)+$signed(-sharing130_r)+$signed(sharing166_r)+$signed(sharing167_r)+$signed(sharing183_r)+$signed(-sharing184_r)+$signed(sharing211_r)+$signed(sharing223_r)+$signed(-sharing224_r)+$signed(sharing233_r)+$signed(sharing244_r)+$signed(0);
assign weighted_sum[19] = $signed(-{in[160],1'b0})+$signed(-in[128])+$signed(in[258])+$signed(-{in[131],1'b0})+$signed({in[451],1'b0})+$signed(-{in[483],1'b0})+$signed({in[452],1'b0})+$signed(-in[133])+$signed(-{in[166],2'b0})+$signed(in[264])+$signed(in[202])+$signed(-{in[395],2'b0})+$signed(-{in[396],2'b0})+$signed(in[268])+$signed(-{in[141],2'b0})+$signed(-in[429])+$signed(-{in[46],1'b0})+$signed(-{in[399],2'b0})+$signed(-in[335])+$signed(in[463])+$signed(-{in[496],1'b0})+$signed(-in[48])+$signed(in[112])+$signed(-in[498])+$signed({in[211],1'b0})+$signed(-in[147])+$signed({in[276],1'b0})+$signed(-in[148])+$signed(in[87])+$signed(-{in[409],2'b0})+$signed(-in[90])+$signed(in[378])+$signed(-in[442])+$signed({in[219],1'b0})+$signed(in[252])+$signed(in[284])+$signed({in[253],1'b0})+$signed(-{in[382],2'b0})+$signed(sharing8_r)+$signed(-sharing9_r)+$signed(sharing54_r)+$signed(sharing55_r)+$signed(sharing86_r)+$signed(sharing87_r)+$signed(sharing118_r)+$signed(sharing119_r)+$signed(sharing143_r)+$signed(sharing144_r)+$signed(sharing168_r)+$signed(sharing187_r)+$signed(-sharing188_r)+$signed(sharing225_r)+$signed(sharing239_r)+$signed(-sharing241_r)+$signed(sharing250_r)+$signed(1);
assign weighted_sum[20] = $signed(-{in[480],1'b0})+$signed(in[449])+$signed({in[34],1'b0})+$signed(-{in[418],1'b0})+$signed({in[323],1'b0})+$signed(-in[3])+$signed(-in[99])+$signed(-in[419])+$signed(-in[68])+$signed(in[356])+$signed(-{in[453],1'b0})+$signed(in[223])+$signed(-in[455])+$signed(-in[7])+$signed(in[167])+$signed({in[424],1'b0})+$signed(-in[40])+$signed(in[233])+$signed(-in[298])+$signed(-in[492])+$signed(-in[301])+$signed(-{in[142],1'b0})+$signed(-in[206])+$signed(-{in[271],1'b0})+$signed(in[241])+$signed(in[497])+$signed(-in[275])+$signed({in[373],1'b0})+$signed(in[21])+$signed({in[310],1'b0})+$signed(-in[282])+$signed(-{in[123],1'b0})+$signed(-in[283])+$signed(in[411])+$signed(in[317])+$signed({in[414],1'b0})+$signed(-in[158])+$signed(in[383])+$signed(sharing22_r)+$signed(-sharing23_r)+$signed(sharing34_r)+$signed(-sharing35_r)+$signed(sharing90_r)+$signed(-sharing91_r)+$signed(sharing122_r)+$signed(-sharing123_r)+$signed(sharing145_r)+$signed(sharing146_r)+$signed(sharing169_r)+$signed(sharing192_r)+$signed(-sharing211_r)+$signed(-sharing219_r)+$signed(sharing237_r)+$signed(sharing240_r)+$signed(-2);
assign weighted_sum[21] = $signed(-in[222])+$signed(in[482])+$signed(-{in[419],1'b0})+$signed(-{in[451],1'b0})+$signed(-in[99])+$signed(-{in[191],1'b0})+$signed({in[356],1'b0})+$signed(-{in[391],2'b0})+$signed(-{in[455],1'b0})+$signed(-in[423])+$signed(in[264])+$signed(-{in[426],2'b0})+$signed({in[492],2'b0})+$signed(-in[300])+$signed(in[269])+$signed(in[45])+$signed({in[334],1'b0})+$signed(in[206])+$signed(in[398])+$signed({in[335],1'b0})+$signed(-in[112])+$signed({in[465],1'b0})+$signed(-in[113])+$signed(in[275])+$signed(in[371])+$signed(-in[405])+$signed(-{in[438],2'b0})+$signed(-{in[406],1'b0})+$signed({in[311],1'b0})+$signed(-{in[439],1'b0})+$signed({in[152],1'b0})+$signed(-{in[442],1'b0})+$signed(-{in[187],1'b0})+$signed(-in[27])+$signed(-in[62])+$signed(in[475])+$signed({in[476],1'b0})+$signed(-in[412])+$signed(in[253])+$signed({in[478],2'b0})+$signed(in[446])+$signed({in[479],2'b0})+$signed({in[95],1'b0})+$signed(sharing26_r)+$signed(sharing27_r)+$signed(sharing62_r)+$signed(-sharing63_r)+$signed(sharing88_r)+$signed(-sharing89_r)+$signed(sharing110_r)+$signed(-sharing111_r)+$signed(sharing136_r)+$signed(-sharing137_r)+$signed(sharing156_r)+$signed(-sharing157_r)+$signed(sharing181_r)+$signed(-sharing182_r)+$signed(sharing201_r)+$signed(sharing229_r)+$signed(sharing246_r)+$signed(2);
assign weighted_sum[22] = $signed({in[384],1'b0})+$signed(in[128])+$signed({in[225],1'b0})+$signed(-in[1])+$signed({in[226],1'b0})+$signed({in[227],2'b0})+$signed(in[451])+$signed({in[100],1'b0})+$signed(in[228])+$signed({in[102],1'b0})+$signed(in[262])+$signed(-in[40])+$signed(-in[73])+$signed(in[490])+$signed({in[44],1'b0})+$signed(-in[12])+$signed(in[140])+$signed({in[397],1'b0})+$signed({in[270],1'b0})+$signed({in[462],1'b0})+$signed({in[463],1'b0})+$signed(-in[79])+$signed(in[271])+$signed(in[112])+$signed({in[113],1'b0})+$signed({in[213],2'b0})+$signed({in[469],1'b0})+$signed({in[214],2'b0})+$signed(in[374])+$signed({in[87],1'b0})+$signed({in[88],1'b0})+$signed({in[57],1'b0})+$signed(-in[409])+$signed(in[441])+$signed(in[473])+$signed(-in[27])+$signed({in[284],1'b0})+$signed(in[124])+$signed(in[477])+$signed({in[127],1'b0})+$signed(sharing10_r)+$signed(-sharing11_r)+$signed(sharing46_r)+$signed(-sharing47_r)+$signed(sharing74_r)+$signed(-sharing75_r)+$signed(sharing96_r)+$signed(-sharing97_r)+$signed(sharing132_r)+$signed(-sharing133_r)+$signed(sharing170_r)+$signed(sharing171_r)+$signed(sharing193_r)+$signed(sharing207_r)+$signed(-sharing208_r)+$signed(0);
assign weighted_sum[23] = $signed({in[256],2'b0})+$signed({in[257],2'b0})+$signed(-in[353])+$signed(-in[193])+$signed(in[33])+$signed(in[162])+$signed(in[418])+$signed(-in[387])+$signed(-{in[388],1'b0})+$signed({in[391],1'b0})+$signed(-in[7])+$signed({in[199],1'b0})+$signed(-in[167])+$signed({in[392],1'b0})+$signed(-in[296])+$signed(-{in[9],1'b0})+$signed({in[73],1'b0})+$signed({in[74],2'b0})+$signed(-in[362])+$signed(in[394])+$signed(in[300])+$signed(-in[205])+$signed({in[238],1'b0})+$signed({in[367],1'b0})+$signed(-in[15])+$signed(-in[399])+$signed(-in[50])+$signed(in[370])+$signed({in[243],2'b0})+$signed(-{in[51],1'b0})+$signed({in[212],2'b0})+$signed(in[117])+$signed(-{in[23],2'b0})+$signed(in[439])+$signed(-in[24])+$signed(-in[59])+$signed(-in[188])+$signed(-in[125])+$signed(in[254])+$signed({in[255],2'b0})+$signed({in[159],1'b0})+$signed(in[127])+$signed(sharing16_r)+$signed(-sharing17_r)+$signed(sharing42_r)+$signed(-sharing43_r)+$signed(sharing64_r)+$signed(-sharing65_r)+$signed(sharing118_r)+$signed(-sharing119_r)+$signed(sharing131_r)+$signed(sharing176_r)+$signed(-sharing193_r)+$signed(-sharing251_r)+$signed(-sharing253_r)+$signed(1);
assign weighted_sum[24] = $signed(-{in[289],1'b0})+$signed(-{in[257],1'b0})+$signed(-in[130])+$signed(in[194])+$signed({in[131],1'b0})+$signed(in[483])+$signed(in[421])+$signed(in[200])+$signed(in[360])+$signed(in[361])+$signed({in[268],1'b0})+$signed(-{in[269],1'b0})+$signed(in[237])+$signed(-{in[270],1'b0})+$signed({in[496],1'b0})+$signed(-in[51])+$signed(in[211])+$signed(in[20])+$signed(in[468])+$signed(-{in[245],2'b0})+$signed(in[437])+$signed(in[406])+$signed(in[375])+$signed(-in[56])+$signed(-{in[441],1'b0})+$signed(in[409])+$signed(-{in[154],2'b0})+$signed(-in[250])+$signed(in[314])+$signed(in[346])+$signed(in[476])+$signed(-in[95])+$signed(sharing28_r)+$signed(sharing29_r)+$signed(sharing56_r)+$signed(sharing57_r)+$signed(sharing88_r)+$signed(sharing89_r)+$signed(sharing120_r)+$signed(sharing121_r)+$signed(sharing147_r)+$signed(sharing148_r)+$signed(sharing172_r)+$signed(sharing194_r)+$signed(sharing195_r)+$signed(sharing212_r)+$signed(sharing213_r)+$signed(sharing226_r)+$signed(sharing234_r)+$signed(sharing239_r)+$signed(sharing245_r)+$signed(sharing251_r)+$signed(2);
assign weighted_sum[25] = $signed({in[254],1'b0})+$signed(-in[0])+$signed({in[34],2'b0})+$signed({in[483],1'b0})+$signed(-in[421])+$signed(-in[165])+$signed(-in[329])+$signed(in[425])+$signed(-in[74])+$signed({in[459],2'b0})+$signed({in[491],1'b0})+$signed({in[460],2'b0})+$signed({in[141],1'b0})+$signed(-{in[430],1'b0})+$signed(in[462])+$signed({in[463],1'b0})+$signed({in[464],1'b0})+$signed({in[145],1'b0})+$signed(in[49])+$signed(in[498])+$signed(in[470])+$signed({in[472],2'b0})+$signed(-in[280])+$signed({in[473],2'b0})+$signed(in[441])+$signed(-{in[316],1'b0})+$signed(in[188])+$signed({in[477],1'b0})+$signed({in[126],1'b0})+$signed({in[415],1'b0})+$signed(-in[159])+$signed(sharing2_r)+$signed(-sharing3_r)+$signed(sharing58_r)+$signed(sharing59_r)+$signed(sharing90_r)+$signed(sharing91_r)+$signed(sharing112_r)+$signed(-sharing113_r)+$signed(sharing141_r)+$signed(-sharing142_r)+$signed(sharing172_r)+$signed(sharing196_r)+$signed(sharing197_r)+$signed(sharing227_r)+$signed(sharing246_r)+$signed(sharing252_r)+$signed(sharing254_r)+$signed(sharing255_r)+$signed(0);
assign weighted_sum[26] = $signed(-in[96])+$signed(-{in[257],1'b0})+$signed(in[95])+$signed(-{in[292],1'b0})+$signed(in[388])+$signed({in[229],1'b0})+$signed(-{in[231],1'b0})+$signed({in[167],1'b0})+$signed(in[319])+$signed({in[361],1'b0})+$signed(in[10])+$signed(in[107])+$signed(in[203])+$signed(in[76])+$signed(in[238])+$signed(-in[463])+$signed(-in[242])+$signed(-{in[243],1'b0})+$signed(-{in[244],1'b0})+$signed(in[500])+$signed(-in[85])+$signed(-{in[406],1'b0})+$signed({in[375],1'b0})+$signed(-in[439])+$signed(-{in[441],2'b0})+$signed(-in[345])+$signed(-in[506])+$signed({in[188],1'b0})+$signed({in[252],1'b0})+$signed({in[412],1'b0})+$signed({in[253],2'b0})+$signed({in[189],1'b0})+$signed(in[93])+$signed({in[444],1'b0})+$signed({in[158],1'b0})+$signed({in[446],1'b0})+$signed(-{in[255],1'b0})+$signed(in[447])+$signed(sharing6_r)+$signed(-sharing7_r)+$signed(sharing58_r)+$signed(-sharing59_r)+$signed(sharing66_r)+$signed(-sharing67_r)+$signed(sharing122_r)+$signed(sharing123_r)+$signed(sharing149_r)+$signed(sharing150_r)+$signed(sharing166_r)+$signed(-sharing167_r)+$signed(sharing198_r)+$signed(sharing214_r)+$signed(sharing215_r)+$signed(sharing228_r)+$signed(sharing235_r)+$signed(3);
assign weighted_sum[27] = $signed({in[448],2'b0})+$signed({in[288],1'b0})+$signed(in[192])+$signed({in[98],1'b0})+$signed(in[99])+$signed({in[388],1'b0})+$signed(in[389])+$signed(-in[261])+$signed({in[38],1'b0})+$signed(-{in[102],1'b0})+$signed(-in[70])+$signed(-in[135])+$signed(in[266])+$signed(in[490])+$signed(in[139])+$signed(in[395])+$signed({in[493],1'b0})+$signed({in[462],1'b0})+$signed({in[207],1'b0})+$signed({in[111],1'b0})+$signed(-in[495])+$signed(-in[144])+$signed(-in[240])+$signed(in[400])+$signed(-{in[210],1'b0})+$signed(-in[274])+$signed({in[436],1'b0})+$signed(in[213])+$signed(-in[405])+$signed(-in[150])+$signed(-in[470])+$signed({in[279],1'b0})+$signed({in[503],1'b0})+$signed({in[504],1'b0})+$signed(in[153])+$signed({in[154],1'b0})+$signed({in[314],1'b0})+$signed(-in[410])+$signed(-{in[442],1'b0})+$signed(-in[252])+$signed(-in[284])+$signed({in[479],1'b0})+$signed(in[415])+$signed(sharing28_r)+$signed(-sharing29_r)+$signed(sharing60_r)+$signed(sharing61_r)+$signed(sharing80_r)+$signed(-sharing81_r)+$signed(sharing124_r)+$signed(sharing125_r)+$signed(sharing173_r)+$signed(sharing216_r)+$signed(sharing247_r)+$signed(0);
assign weighted_sum[28] = $signed(-{in[64],2'b0})+$signed(in[257])+$signed(-in[225])+$signed(in[162])+$signed(in[354])+$signed(in[323])+$signed(in[419])+$signed(in[483])+$signed({in[228],1'b0})+$signed(in[324])+$signed(-{in[389],2'b0})+$signed(in[198])+$signed({in[46],2'b0})+$signed({in[47],1'b0})+$signed(-in[239])+$signed(-in[303])+$signed(in[80])+$signed(-{in[402],2'b0})+$signed(in[466])+$signed(-{in[51],2'b0})+$signed({in[467],1'b0})+$signed(-in[243])+$signed(in[404])+$signed(in[405])+$signed(-in[438])+$signed(-in[23])+$signed({in[216],1'b0})+$signed(in[216])+$signed({in[408],1'b0})+$signed({in[409],1'b0})+$signed(in[473])+$signed(-{in[379],1'b0})+$signed(-{in[380],1'b0})+$signed(-in[413])+$signed({in[254],1'b0})+$signed(-in[414])+$signed(sharing20_r)+$signed(-sharing21_r)+$signed(sharing40_r)+$signed(-sharing41_r)+$signed(sharing92_r)+$signed(sharing93_r)+$signed(sharing126_r)+$signed(sharing149_r)+$signed(-sharing150_r)+$signed(-sharing168_r)+$signed(sharing199_r)+$signed(sharing200_r)+$signed(sharing202_r)+$signed(sharing229_r)+$signed(sharing242_r)+$signed(1);
assign weighted_sum[29] = $signed(-in[384])+$signed(in[192])+$signed(in[416])+$signed(in[450])+$signed(in[290])+$signed(-{in[131],2'b0})+$signed({in[67],1'b0})+$signed(in[131])+$signed({in[419],2'b0})+$signed(in[419])+$signed({in[388],1'b0})+$signed({in[420],2'b0})+$signed({in[69],2'b0})+$signed({in[389],1'b0})+$signed({in[70],3'b0})+$signed(in[487])+$signed(-in[74])+$signed(in[298])+$signed(-in[491])+$signed(-{in[397],1'b0})+$signed(-in[301])+$signed(in[365])+$signed({in[430],1'b0})+$signed({in[240],2'b0})+$signed(-in[368])+$signed({in[81],2'b0})+$signed({in[241],1'b0})+$signed(in[241])+$signed(-in[146])+$signed(-{in[19],1'b0})+$signed(-{in[468],1'b0})+$signed(-{in[21],1'b0})+$signed(-in[213])+$signed(-in[118])+$signed(-in[54])+$signed(in[248])+$signed({in[409],2'b0})+$signed(-{in[506],1'b0})+$signed({in[251],2'b0})+$signed(-in[219])+$signed(in[284])+$signed(sharing14_r)+$signed(-sharing15_r)+$signed(sharing62_r)+$signed(sharing63_r)+$signed(sharing68_r)+$signed(-sharing69_r)+$signed(sharing120_r)+$signed(-sharing121_r)+$signed(sharing151_r)+$signed(sharing152_r)+$signed(sharing174_r)+$signed(sharing175_r)+$signed(-sharing203_r)+$signed(sharing228_r)+$signed(-sharing230_r)+$signed(2);
assign weighted_sum[30] = $signed(-in[128])+$signed(-{in[193],1'b0})+$signed(-in[129])+$signed({in[258],1'b0})+$signed(-in[162])+$signed(-in[322])+$signed(-{in[387],2'b0})+$signed(-{in[37],1'b0})+$signed(-{in[421],1'b0})+$signed({in[262],1'b0})+$signed(-in[70])+$signed({in[327],1'b0})+$signed({in[328],1'b0})+$signed(-{in[233],1'b0})+$signed(-{in[425],1'b0})+$signed({in[236],1'b0})+$signed(-in[204])+$signed(-{in[428],1'b0})+$signed({in[237],1'b0})+$signed(-{in[493],1'b0})+$signed(-in[334])+$signed(-in[398])+$signed(-{in[399],1'b0})+$signed(-{in[400],2'b0})+$signed(-{in[304],1'b0})+$signed(-{in[401],2'b0})+$signed(-in[82])+$signed(-{in[51],1'b0})+$signed({in[53],1'b0})+$signed({in[405],1'b0})+$signed(-{in[246],2'b0})+$signed(in[54])+$signed(-in[502])+$signed(-{in[24],2'b0})+$signed(-{in[216],1'b0})+$signed(-{in[280],1'b0})+$signed(in[441])+$signed(-in[154])+$signed({in[251],1'b0})+$signed(in[27])+$signed(-in[475])+$signed(-{in[220],1'b0})+$signed(in[60])+$signed(-{in[414],2'b0})+$signed(-{in[415],2'b0})+$signed(in[383])+$signed(sharing30_r)+$signed(sharing31_r)+$signed(sharing52_r)+$signed(-sharing53_r)+$signed(sharing94_r)+$signed(sharing95_r)+$signed(sharing114_r)+$signed(-sharing115_r)+$signed(sharing153_r)+$signed(sharing154_r)+$signed(-sharing169_r)+$signed(sharing178_r)+$signed(-sharing179_r)+$signed(sharing214_r)+$signed(-sharing215_r)+$signed(-sharing227_r)+$signed(1);
assign weighted_sum[31] = $signed(-in[258])+$signed(-in[418])+$signed({in[483],1'b0})+$signed(-{in[387],1'b0})+$signed(-in[35])+$signed(in[388])+$signed({in[229],1'b0})+$signed({in[293],1'b0})+$signed({in[230],2'b0})+$signed(-in[38])+$signed({in[231],2'b0})+$signed({in[232],1'b0})+$signed(in[456])+$signed(in[330])+$signed(-in[75])+$signed(-{in[76],1'b0})+$signed(in[237])+$signed(in[333])+$signed(-in[493])+$signed({in[111],1'b0})+$signed(-in[175])+$signed({in[144],1'b0})+$signed(in[48])+$signed({in[368],1'b0})+$signed({in[241],2'b0})+$signed(in[244])+$signed(in[469])+$signed(-in[55])+$signed(in[471])+$signed(-{in[24],1'b0})+$signed(-in[88])+$signed({in[281],1'b0})+$signed(-in[89])+$signed({in[59],1'b0})+$signed(in[59])+$signed(in[123])+$signed({in[60],2'b0})+$signed({in[28],1'b0})+$signed(-in[155])+$signed(-{in[413],1'b0})+$signed(in[317])+$signed({in[62],1'b0})+$signed(in[318])+$signed({in[63],1'b0})+$signed(sharing30_r)+$signed(-sharing31_r)+$signed(sharing44_r)+$signed(-sharing45_r)+$signed(sharing84_r)+$signed(-sharing85_r)+$signed(sharing102_r)+$signed(-sharing103_r)+$signed(sharing151_r)+$signed(-sharing152_r)+$signed(sharing176_r)+$signed(-sharing198_r)+$signed(2);
assign out[0] = (weighted_sum[0][9]==1) ? 4'd0 : (weighted_sum[0][8:2] > 6 ? 4'd6 : weighted_sum[0][5:2]);
assign out[1] = (weighted_sum[1][9]==1) ? 4'd0 : (weighted_sum[1][8:2] > 6 ? 4'd6 : weighted_sum[1][5:2]);
assign out[2] = (weighted_sum[2][9]==1) ? 4'd0 : (weighted_sum[2][8:2] > 6 ? 4'd6 : weighted_sum[2][5:2]);
assign out[3] = (weighted_sum[3][9]==1) ? 4'd0 : (weighted_sum[3][8:2] > 6 ? 4'd6 : weighted_sum[3][5:2]);
assign out[4] = (weighted_sum[4][9]==1) ? 4'd0 : (weighted_sum[4][8:2] > 6 ? 4'd6 : weighted_sum[4][5:2]);
assign out[5] = (weighted_sum[5][9]==1) ? 4'd0 : (weighted_sum[5][8:2] > 6 ? 4'd6 : weighted_sum[5][5:2]);
assign out[6] = (weighted_sum[6][9]==1) ? 4'd0 : (weighted_sum[6][8:2] > 6 ? 4'd6 : weighted_sum[6][5:2]);
assign out[7] = (weighted_sum[7][9]==1) ? 4'd0 : (weighted_sum[7][8:2] > 6 ? 4'd6 : weighted_sum[7][5:2]);
assign out[8] = (weighted_sum[8][9]==1) ? 4'd0 : (weighted_sum[8][8:2] > 6 ? 4'd6 : weighted_sum[8][5:2]);
assign out[9] = (weighted_sum[9][9]==1) ? 4'd0 : (weighted_sum[9][8:2] > 6 ? 4'd6 : weighted_sum[9][5:2]);
assign out[10] = (weighted_sum[10][9]==1) ? 4'd0 : (weighted_sum[10][8:2] > 6 ? 4'd6 : weighted_sum[10][5:2]);
assign out[11] = (weighted_sum[11][9]==1) ? 4'd0 : (weighted_sum[11][8:2] > 6 ? 4'd6 : weighted_sum[11][5:2]);
assign out[12] = (weighted_sum[12][9]==1) ? 4'd0 : (weighted_sum[12][8:2] > 6 ? 4'd6 : weighted_sum[12][5:2]);
assign out[13] = (weighted_sum[13][9]==1) ? 4'd0 : (weighted_sum[13][8:2] > 6 ? 4'd6 : weighted_sum[13][5:2]);
assign out[14] = (weighted_sum[14][9]==1) ? 4'd0 : (weighted_sum[14][8:2] > 6 ? 4'd6 : weighted_sum[14][5:2]);
assign out[15] = (weighted_sum[15][9]==1) ? 4'd0 : (weighted_sum[15][8:2] > 6 ? 4'd6 : weighted_sum[15][5:2]);
assign out[16] = (weighted_sum[16][9]==1) ? 4'd0 : (weighted_sum[16][8:2] > 6 ? 4'd6 : weighted_sum[16][5:2]);
assign out[17] = (weighted_sum[17][9]==1) ? 4'd0 : (weighted_sum[17][8:2] > 6 ? 4'd6 : weighted_sum[17][5:2]);
assign out[18] = (weighted_sum[18][9]==1) ? 4'd0 : (weighted_sum[18][8:2] > 6 ? 4'd6 : weighted_sum[18][5:2]);
assign out[19] = (weighted_sum[19][9]==1) ? 4'd0 : (weighted_sum[19][8:2] > 6 ? 4'd6 : weighted_sum[19][5:2]);
assign out[20] = (weighted_sum[20][9]==1) ? 4'd0 : (weighted_sum[20][8:2] > 6 ? 4'd6 : weighted_sum[20][5:2]);
assign out[21] = (weighted_sum[21][9]==1) ? 4'd0 : (weighted_sum[21][8:2] > 6 ? 4'd6 : weighted_sum[21][5:2]);
assign out[22] = (weighted_sum[22][9]==1) ? 4'd0 : (weighted_sum[22][8:2] > 6 ? 4'd6 : weighted_sum[22][5:2]);
assign out[23] = (weighted_sum[23][9]==1) ? 4'd0 : (weighted_sum[23][8:2] > 6 ? 4'd6 : weighted_sum[23][5:2]);
assign out[24] = (weighted_sum[24][9]==1) ? 4'd0 : (weighted_sum[24][8:2] > 6 ? 4'd6 : weighted_sum[24][5:2]);
assign out[25] = (weighted_sum[25][9]==1) ? 4'd0 : (weighted_sum[25][8:2] > 6 ? 4'd6 : weighted_sum[25][5:2]);
assign out[26] = (weighted_sum[26][9]==1) ? 4'd0 : (weighted_sum[26][8:2] > 6 ? 4'd6 : weighted_sum[26][5:2]);
assign out[27] = (weighted_sum[27][9]==1) ? 4'd0 : (weighted_sum[27][8:2] > 6 ? 4'd6 : weighted_sum[27][5:2]);
assign out[28] = (weighted_sum[28][9]==1) ? 4'd0 : (weighted_sum[28][8:2] > 6 ? 4'd6 : weighted_sum[28][5:2]);
assign out[29] = (weighted_sum[29][9]==1) ? 4'd0 : (weighted_sum[29][8:2] > 6 ? 4'd6 : weighted_sum[29][5:2]);
assign out[30] = (weighted_sum[30][9]==1) ? 4'd0 : (weighted_sum[30][8:2] > 6 ? 4'd6 : weighted_sum[30][5:2]);
assign out[31] = (weighted_sum[31][9]==1) ? 4'd0 : (weighted_sum[31][8:2] > 6 ? 4'd6 : weighted_sum[31][5:2]);

always_ff @ (posedge clk or posedge rst) begin
	if (rst) begin
		sharing0_r <= 0;
		sharing1_r <= 0;
		sharing2_r <= 0;
		sharing3_r <= 0;
		sharing4_r <= 0;
		sharing5_r <= 0;
		sharing6_r <= 0;
		sharing7_r <= 0;
		sharing8_r <= 0;
		sharing9_r <= 0;
		sharing10_r <= 0;
		sharing11_r <= 0;
		sharing12_r <= 0;
		sharing13_r <= 0;
		sharing14_r <= 0;
		sharing15_r <= 0;
		sharing16_r <= 0;
		sharing17_r <= 0;
		sharing18_r <= 0;
		sharing19_r <= 0;
		sharing20_r <= 0;
		sharing21_r <= 0;
		sharing22_r <= 0;
		sharing23_r <= 0;
		sharing24_r <= 0;
		sharing25_r <= 0;
		sharing26_r <= 0;
		sharing27_r <= 0;
		sharing28_r <= 0;
		sharing29_r <= 0;
		sharing30_r <= 0;
		sharing31_r <= 0;
		sharing32_r <= 0;
		sharing33_r <= 0;
		sharing34_r <= 0;
		sharing35_r <= 0;
		sharing36_r <= 0;
		sharing37_r <= 0;
		sharing38_r <= 0;
		sharing39_r <= 0;
		sharing40_r <= 0;
		sharing41_r <= 0;
		sharing42_r <= 0;
		sharing43_r <= 0;
		sharing44_r <= 0;
		sharing45_r <= 0;
		sharing46_r <= 0;
		sharing47_r <= 0;
		sharing48_r <= 0;
		sharing49_r <= 0;
		sharing50_r <= 0;
		sharing51_r <= 0;
		sharing52_r <= 0;
		sharing53_r <= 0;
		sharing54_r <= 0;
		sharing55_r <= 0;
		sharing56_r <= 0;
		sharing57_r <= 0;
		sharing58_r <= 0;
		sharing59_r <= 0;
		sharing60_r <= 0;
		sharing61_r <= 0;
		sharing62_r <= 0;
		sharing63_r <= 0;
		sharing64_r <= 0;
		sharing65_r <= 0;
		sharing66_r <= 0;
		sharing67_r <= 0;
		sharing68_r <= 0;
		sharing69_r <= 0;
		sharing70_r <= 0;
		sharing71_r <= 0;
		sharing72_r <= 0;
		sharing73_r <= 0;
		sharing74_r <= 0;
		sharing75_r <= 0;
		sharing76_r <= 0;
		sharing77_r <= 0;
		sharing78_r <= 0;
		sharing79_r <= 0;
		sharing80_r <= 0;
		sharing81_r <= 0;
		sharing82_r <= 0;
		sharing83_r <= 0;
		sharing84_r <= 0;
		sharing85_r <= 0;
		sharing86_r <= 0;
		sharing87_r <= 0;
		sharing88_r <= 0;
		sharing89_r <= 0;
		sharing90_r <= 0;
		sharing91_r <= 0;
		sharing92_r <= 0;
		sharing93_r <= 0;
		sharing94_r <= 0;
		sharing95_r <= 0;
		sharing96_r <= 0;
		sharing97_r <= 0;
		sharing98_r <= 0;
		sharing99_r <= 0;
		sharing100_r <= 0;
		sharing101_r <= 0;
		sharing102_r <= 0;
		sharing103_r <= 0;
		sharing104_r <= 0;
		sharing105_r <= 0;
		sharing106_r <= 0;
		sharing107_r <= 0;
		sharing108_r <= 0;
		sharing109_r <= 0;
		sharing110_r <= 0;
		sharing111_r <= 0;
		sharing112_r <= 0;
		sharing113_r <= 0;
		sharing114_r <= 0;
		sharing115_r <= 0;
		sharing116_r <= 0;
		sharing117_r <= 0;
		sharing118_r <= 0;
		sharing119_r <= 0;
		sharing120_r <= 0;
		sharing121_r <= 0;
		sharing122_r <= 0;
		sharing123_r <= 0;
		sharing124_r <= 0;
		sharing125_r <= 0;
		sharing126_r <= 0;
		sharing127_r <= 0;
		sharing128_r <= 0;
		sharing129_r <= 0;
		sharing130_r <= 0;
		sharing131_r <= 0;
		sharing132_r <= 0;
		sharing133_r <= 0;
		sharing134_r <= 0;
		sharing135_r <= 0;
		sharing136_r <= 0;
		sharing137_r <= 0;
		sharing138_r <= 0;
		sharing139_r <= 0;
		sharing140_r <= 0;
		sharing141_r <= 0;
		sharing142_r <= 0;
		sharing143_r <= 0;
		sharing144_r <= 0;
		sharing145_r <= 0;
		sharing146_r <= 0;
		sharing147_r <= 0;
		sharing148_r <= 0;
		sharing149_r <= 0;
		sharing150_r <= 0;
		sharing151_r <= 0;
		sharing152_r <= 0;
		sharing153_r <= 0;
		sharing154_r <= 0;
		sharing155_r <= 0;
		sharing156_r <= 0;
		sharing157_r <= 0;
		sharing158_r <= 0;
		sharing159_r <= 0;
		sharing160_r <= 0;
		sharing161_r <= 0;
		sharing162_r <= 0;
		sharing163_r <= 0;
		sharing164_r <= 0;
		sharing165_r <= 0;
		sharing166_r <= 0;
		sharing167_r <= 0;
		sharing168_r <= 0;
		sharing169_r <= 0;
		sharing170_r <= 0;
		sharing171_r <= 0;
		sharing172_r <= 0;
		sharing173_r <= 0;
		sharing174_r <= 0;
		sharing175_r <= 0;
		sharing176_r <= 0;
		sharing177_r <= 0;
		sharing178_r <= 0;
		sharing179_r <= 0;
		sharing180_r <= 0;
		sharing181_r <= 0;
		sharing182_r <= 0;
		sharing183_r <= 0;
		sharing184_r <= 0;
		sharing185_r <= 0;
		sharing186_r <= 0;
		sharing187_r <= 0;
		sharing188_r <= 0;
		sharing189_r <= 0;
		sharing190_r <= 0;
		sharing191_r <= 0;
		sharing192_r <= 0;
		sharing193_r <= 0;
		sharing194_r <= 0;
		sharing195_r <= 0;
		sharing196_r <= 0;
		sharing197_r <= 0;
		sharing198_r <= 0;
		sharing199_r <= 0;
		sharing200_r <= 0;
		sharing201_r <= 0;
		sharing202_r <= 0;
		sharing203_r <= 0;
		sharing204_r <= 0;
		sharing205_r <= 0;
		sharing206_r <= 0;
		sharing207_r <= 0;
		sharing208_r <= 0;
		sharing209_r <= 0;
		sharing210_r <= 0;
		sharing211_r <= 0;
		sharing212_r <= 0;
		sharing213_r <= 0;
		sharing214_r <= 0;
		sharing215_r <= 0;
		sharing216_r <= 0;
		sharing217_r <= 0;
		sharing218_r <= 0;
		sharing219_r <= 0;
		sharing220_r <= 0;
		sharing221_r <= 0;
		sharing222_r <= 0;
		sharing223_r <= 0;
		sharing224_r <= 0;
		sharing225_r <= 0;
		sharing226_r <= 0;
		sharing227_r <= 0;
		sharing228_r <= 0;
		sharing229_r <= 0;
		sharing230_r <= 0;
		sharing231_r <= 0;
		sharing232_r <= 0;
		sharing233_r <= 0;
		sharing234_r <= 0;
		sharing235_r <= 0;
		sharing236_r <= 0;
		sharing237_r <= 0;
		sharing238_r <= 0;
		sharing239_r <= 0;
		sharing240_r <= 0;
		sharing241_r <= 0;
		sharing242_r <= 0;
		sharing243_r <= 0;
		sharing244_r <= 0;
		sharing245_r <= 0;
		sharing246_r <= 0;
		sharing247_r <= 0;
		sharing248_r <= 0;
		sharing249_r <= 0;
		sharing250_r <= 0;
		sharing251_r <= 0;
		sharing252_r <= 0;
		sharing253_r <= 0;
		sharing254_r <= 0;
		sharing255_r <= 0;
	end
	else begin
		sharing0_r <= sharing0_w;
		sharing1_r <= sharing1_w;
		sharing2_r <= sharing2_w;
		sharing3_r <= sharing3_w;
		sharing4_r <= sharing4_w;
		sharing5_r <= sharing5_w;
		sharing6_r <= sharing6_w;
		sharing7_r <= sharing7_w;
		sharing8_r <= sharing8_w;
		sharing9_r <= sharing9_w;
		sharing10_r <= sharing10_w;
		sharing11_r <= sharing11_w;
		sharing12_r <= sharing12_w;
		sharing13_r <= sharing13_w;
		sharing14_r <= sharing14_w;
		sharing15_r <= sharing15_w;
		sharing16_r <= sharing16_w;
		sharing17_r <= sharing17_w;
		sharing18_r <= sharing18_w;
		sharing19_r <= sharing19_w;
		sharing20_r <= sharing20_w;
		sharing21_r <= sharing21_w;
		sharing22_r <= sharing22_w;
		sharing23_r <= sharing23_w;
		sharing24_r <= sharing24_w;
		sharing25_r <= sharing25_w;
		sharing26_r <= sharing26_w;
		sharing27_r <= sharing27_w;
		sharing28_r <= sharing28_w;
		sharing29_r <= sharing29_w;
		sharing30_r <= sharing30_w;
		sharing31_r <= sharing31_w;
		sharing32_r <= sharing32_w;
		sharing33_r <= sharing33_w;
		sharing34_r <= sharing34_w;
		sharing35_r <= sharing35_w;
		sharing36_r <= sharing36_w;
		sharing37_r <= sharing37_w;
		sharing38_r <= sharing38_w;
		sharing39_r <= sharing39_w;
		sharing40_r <= sharing40_w;
		sharing41_r <= sharing41_w;
		sharing42_r <= sharing42_w;
		sharing43_r <= sharing43_w;
		sharing44_r <= sharing44_w;
		sharing45_r <= sharing45_w;
		sharing46_r <= sharing46_w;
		sharing47_r <= sharing47_w;
		sharing48_r <= sharing48_w;
		sharing49_r <= sharing49_w;
		sharing50_r <= sharing50_w;
		sharing51_r <= sharing51_w;
		sharing52_r <= sharing52_w;
		sharing53_r <= sharing53_w;
		sharing54_r <= sharing54_w;
		sharing55_r <= sharing55_w;
		sharing56_r <= sharing56_w;
		sharing57_r <= sharing57_w;
		sharing58_r <= sharing58_w;
		sharing59_r <= sharing59_w;
		sharing60_r <= sharing60_w;
		sharing61_r <= sharing61_w;
		sharing62_r <= sharing62_w;
		sharing63_r <= sharing63_w;
		sharing64_r <= sharing64_w;
		sharing65_r <= sharing65_w;
		sharing66_r <= sharing66_w;
		sharing67_r <= sharing67_w;
		sharing68_r <= sharing68_w;
		sharing69_r <= sharing69_w;
		sharing70_r <= sharing70_w;
		sharing71_r <= sharing71_w;
		sharing72_r <= sharing72_w;
		sharing73_r <= sharing73_w;
		sharing74_r <= sharing74_w;
		sharing75_r <= sharing75_w;
		sharing76_r <= sharing76_w;
		sharing77_r <= sharing77_w;
		sharing78_r <= sharing78_w;
		sharing79_r <= sharing79_w;
		sharing80_r <= sharing80_w;
		sharing81_r <= sharing81_w;
		sharing82_r <= sharing82_w;
		sharing83_r <= sharing83_w;
		sharing84_r <= sharing84_w;
		sharing85_r <= sharing85_w;
		sharing86_r <= sharing86_w;
		sharing87_r <= sharing87_w;
		sharing88_r <= sharing88_w;
		sharing89_r <= sharing89_w;
		sharing90_r <= sharing90_w;
		sharing91_r <= sharing91_w;
		sharing92_r <= sharing92_w;
		sharing93_r <= sharing93_w;
		sharing94_r <= sharing94_w;
		sharing95_r <= sharing95_w;
		sharing96_r <= sharing96_w;
		sharing97_r <= sharing97_w;
		sharing98_r <= sharing98_w;
		sharing99_r <= sharing99_w;
		sharing100_r <= sharing100_w;
		sharing101_r <= sharing101_w;
		sharing102_r <= sharing102_w;
		sharing103_r <= sharing103_w;
		sharing104_r <= sharing104_w;
		sharing105_r <= sharing105_w;
		sharing106_r <= sharing106_w;
		sharing107_r <= sharing107_w;
		sharing108_r <= sharing108_w;
		sharing109_r <= sharing109_w;
		sharing110_r <= sharing110_w;
		sharing111_r <= sharing111_w;
		sharing112_r <= sharing112_w;
		sharing113_r <= sharing113_w;
		sharing114_r <= sharing114_w;
		sharing115_r <= sharing115_w;
		sharing116_r <= sharing116_w;
		sharing117_r <= sharing117_w;
		sharing118_r <= sharing118_w;
		sharing119_r <= sharing119_w;
		sharing120_r <= sharing120_w;
		sharing121_r <= sharing121_w;
		sharing122_r <= sharing122_w;
		sharing123_r <= sharing123_w;
		sharing124_r <= sharing124_w;
		sharing125_r <= sharing125_w;
		sharing126_r <= sharing126_w;
		sharing127_r <= sharing127_w;
		sharing128_r <= sharing128_w;
		sharing129_r <= sharing129_w;
		sharing130_r <= sharing130_w;
		sharing131_r <= sharing131_w;
		sharing132_r <= sharing132_w;
		sharing133_r <= sharing133_w;
		sharing134_r <= sharing134_w;
		sharing135_r <= sharing135_w;
		sharing136_r <= sharing136_w;
		sharing137_r <= sharing137_w;
		sharing138_r <= sharing138_w;
		sharing139_r <= sharing139_w;
		sharing140_r <= sharing140_w;
		sharing141_r <= sharing141_w;
		sharing142_r <= sharing142_w;
		sharing143_r <= sharing143_w;
		sharing144_r <= sharing144_w;
		sharing145_r <= sharing145_w;
		sharing146_r <= sharing146_w;
		sharing147_r <= sharing147_w;
		sharing148_r <= sharing148_w;
		sharing149_r <= sharing149_w;
		sharing150_r <= sharing150_w;
		sharing151_r <= sharing151_w;
		sharing152_r <= sharing152_w;
		sharing153_r <= sharing153_w;
		sharing154_r <= sharing154_w;
		sharing155_r <= sharing155_w;
		sharing156_r <= sharing156_w;
		sharing157_r <= sharing157_w;
		sharing158_r <= sharing158_w;
		sharing159_r <= sharing159_w;
		sharing160_r <= sharing160_w;
		sharing161_r <= sharing161_w;
		sharing162_r <= sharing162_w;
		sharing163_r <= sharing163_w;
		sharing164_r <= sharing164_w;
		sharing165_r <= sharing165_w;
		sharing166_r <= sharing166_w;
		sharing167_r <= sharing167_w;
		sharing168_r <= sharing168_w;
		sharing169_r <= sharing169_w;
		sharing170_r <= sharing170_w;
		sharing171_r <= sharing171_w;
		sharing172_r <= sharing172_w;
		sharing173_r <= sharing173_w;
		sharing174_r <= sharing174_w;
		sharing175_r <= sharing175_w;
		sharing176_r <= sharing176_w;
		sharing177_r <= sharing177_w;
		sharing178_r <= sharing178_w;
		sharing179_r <= sharing179_w;
		sharing180_r <= sharing180_w;
		sharing181_r <= sharing181_w;
		sharing182_r <= sharing182_w;
		sharing183_r <= sharing183_w;
		sharing184_r <= sharing184_w;
		sharing185_r <= sharing185_w;
		sharing186_r <= sharing186_w;
		sharing187_r <= sharing187_w;
		sharing188_r <= sharing188_w;
		sharing189_r <= sharing189_w;
		sharing190_r <= sharing190_w;
		sharing191_r <= sharing191_w;
		sharing192_r <= sharing192_w;
		sharing193_r <= sharing193_w;
		sharing194_r <= sharing194_w;
		sharing195_r <= sharing195_w;
		sharing196_r <= sharing196_w;
		sharing197_r <= sharing197_w;
		sharing198_r <= sharing198_w;
		sharing199_r <= sharing199_w;
		sharing200_r <= sharing200_w;
		sharing201_r <= sharing201_w;
		sharing202_r <= sharing202_w;
		sharing203_r <= sharing203_w;
		sharing204_r <= sharing204_w;
		sharing205_r <= sharing205_w;
		sharing206_r <= sharing206_w;
		sharing207_r <= sharing207_w;
		sharing208_r <= sharing208_w;
		sharing209_r <= sharing209_w;
		sharing210_r <= sharing210_w;
		sharing211_r <= sharing211_w;
		sharing212_r <= sharing212_w;
		sharing213_r <= sharing213_w;
		sharing214_r <= sharing214_w;
		sharing215_r <= sharing215_w;
		sharing216_r <= sharing216_w;
		sharing217_r <= sharing217_w;
		sharing218_r <= sharing218_w;
		sharing219_r <= sharing219_w;
		sharing220_r <= sharing220_w;
		sharing221_r <= sharing221_w;
		sharing222_r <= sharing222_w;
		sharing223_r <= sharing223_w;
		sharing224_r <= sharing224_w;
		sharing225_r <= sharing225_w;
		sharing226_r <= sharing226_w;
		sharing227_r <= sharing227_w;
		sharing228_r <= sharing228_w;
		sharing229_r <= sharing229_w;
		sharing230_r <= sharing230_w;
		sharing231_r <= sharing231_w;
		sharing232_r <= sharing232_w;
		sharing233_r <= sharing233_w;
		sharing234_r <= sharing234_w;
		sharing235_r <= sharing235_w;
		sharing236_r <= sharing236_w;
		sharing237_r <= sharing237_w;
		sharing238_r <= sharing238_w;
		sharing239_r <= sharing239_w;
		sharing240_r <= sharing240_w;
		sharing241_r <= sharing241_w;
		sharing242_r <= sharing242_w;
		sharing243_r <= sharing243_w;
		sharing244_r <= sharing244_w;
		sharing245_r <= sharing245_w;
		sharing246_r <= sharing246_w;
		sharing247_r <= sharing247_w;
		sharing248_r <= sharing248_w;
		sharing249_r <= sharing249_w;
		sharing250_r <= sharing250_w;
		sharing251_r <= sharing251_w;
		sharing252_r <= sharing252_w;
		sharing253_r <= sharing253_w;
		sharing254_r <= sharing254_w;
		sharing255_r <= sharing255_w;
	end
end
endmodule
