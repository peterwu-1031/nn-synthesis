module conv1 (
	input [7:0] in [0:783],
	input clk,
	input rst,
	output [3:0] out [0:506]
);

logic [12:0] weighted_sum [0:506];
logic [12:0] sharing0_r, sharing0_w;
logic [12:0] sharing1_r, sharing1_w;
logic [12:0] sharing2_r, sharing2_w;
logic [12:0] sharing3_r, sharing3_w;
logic [12:0] sharing4_r, sharing4_w;
logic [12:0] sharing5_r, sharing5_w;
logic [12:0] sharing6_r, sharing6_w;
logic [12:0] sharing7_r, sharing7_w;
logic [12:0] sharing8_r, sharing8_w;
logic [12:0] sharing9_r, sharing9_w;
logic [12:0] sharing10_r, sharing10_w;
logic [12:0] sharing11_r, sharing11_w;
logic [12:0] sharing12_r, sharing12_w;
logic [12:0] sharing13_r, sharing13_w;
logic [12:0] sharing14_r, sharing14_w;
logic [12:0] sharing15_r, sharing15_w;
logic [12:0] sharing16_r, sharing16_w;
logic [12:0] sharing17_r, sharing17_w;
logic [12:0] sharing18_r, sharing18_w;
logic [12:0] sharing19_r, sharing19_w;
logic [12:0] sharing20_r, sharing20_w;
logic [12:0] sharing21_r, sharing21_w;
logic [12:0] sharing22_r, sharing22_w;
logic [12:0] sharing23_r, sharing23_w;
logic [12:0] sharing24_r, sharing24_w;
logic [12:0] sharing25_r, sharing25_w;
logic [12:0] sharing26_r, sharing26_w;
logic [12:0] sharing27_r, sharing27_w;
logic [12:0] sharing28_r, sharing28_w;
logic [12:0] sharing29_r, sharing29_w;
logic [12:0] sharing30_r, sharing30_w;
logic [12:0] sharing31_r, sharing31_w;
logic [12:0] sharing32_r, sharing32_w;
logic [12:0] sharing33_r, sharing33_w;
logic [12:0] sharing34_r, sharing34_w;
logic [12:0] sharing35_r, sharing35_w;
logic [12:0] sharing36_r, sharing36_w;
logic [12:0] sharing37_r, sharing37_w;
logic [12:0] sharing38_r, sharing38_w;
logic [12:0] sharing39_r, sharing39_w;
logic [12:0] sharing40_r, sharing40_w;
logic [12:0] sharing41_r, sharing41_w;
logic [12:0] sharing42_r, sharing42_w;
logic [12:0] sharing43_r, sharing43_w;
logic [12:0] sharing44_r, sharing44_w;
logic [12:0] sharing45_r, sharing45_w;
logic [12:0] sharing46_r, sharing46_w;
logic [12:0] sharing47_r, sharing47_w;
logic [12:0] sharing48_r, sharing48_w;
logic [12:0] sharing49_r, sharing49_w;
logic [12:0] sharing50_r, sharing50_w;
logic [12:0] sharing51_r, sharing51_w;
logic [12:0] sharing52_r, sharing52_w;
logic [12:0] sharing53_r, sharing53_w;
logic [12:0] sharing54_r, sharing54_w;
logic [12:0] sharing55_r, sharing55_w;
logic [12:0] sharing56_r, sharing56_w;
logic [12:0] sharing57_r, sharing57_w;
logic [12:0] sharing58_r, sharing58_w;
logic [12:0] sharing59_r, sharing59_w;
logic [12:0] sharing60_r, sharing60_w;
logic [12:0] sharing61_r, sharing61_w;
logic [12:0] sharing62_r, sharing62_w;
logic [12:0] sharing63_r, sharing63_w;
logic [12:0] sharing64_r, sharing64_w;
logic [12:0] sharing65_r, sharing65_w;
logic [12:0] sharing66_r, sharing66_w;
logic [12:0] sharing67_r, sharing67_w;
logic [12:0] sharing68_r, sharing68_w;
logic [12:0] sharing69_r, sharing69_w;
logic [12:0] sharing70_r, sharing70_w;
logic [12:0] sharing71_r, sharing71_w;
logic [12:0] sharing72_r, sharing72_w;
logic [12:0] sharing73_r, sharing73_w;
logic [12:0] sharing74_r, sharing74_w;
logic [12:0] sharing75_r, sharing75_w;
logic [12:0] sharing76_r, sharing76_w;
logic [12:0] sharing77_r, sharing77_w;
logic [12:0] sharing78_r, sharing78_w;
logic [12:0] sharing79_r, sharing79_w;
logic [12:0] sharing80_r, sharing80_w;
logic [12:0] sharing81_r, sharing81_w;
logic [12:0] sharing82_r, sharing82_w;
logic [12:0] sharing83_r, sharing83_w;
logic [12:0] sharing84_r, sharing84_w;
logic [12:0] sharing85_r, sharing85_w;
logic [12:0] sharing86_r, sharing86_w;
logic [12:0] sharing87_r, sharing87_w;
logic [12:0] sharing88_r, sharing88_w;
logic [12:0] sharing89_r, sharing89_w;
logic [12:0] sharing90_r, sharing90_w;
logic [12:0] sharing91_r, sharing91_w;
logic [12:0] sharing92_r, sharing92_w;
logic [12:0] sharing93_r, sharing93_w;
logic [12:0] sharing94_r, sharing94_w;
logic [12:0] sharing95_r, sharing95_w;
logic [12:0] sharing96_r, sharing96_w;
logic [12:0] sharing97_r, sharing97_w;
logic [12:0] sharing98_r, sharing98_w;
logic [12:0] sharing99_r, sharing99_w;
logic [12:0] sharing100_r, sharing100_w;
logic [12:0] sharing101_r, sharing101_w;
logic [12:0] sharing102_r, sharing102_w;
logic [12:0] sharing103_r, sharing103_w;
logic [12:0] sharing104_r, sharing104_w;
logic [12:0] sharing105_r, sharing105_w;
logic [12:0] sharing106_r, sharing106_w;
logic [12:0] sharing107_r, sharing107_w;
logic [12:0] sharing108_r, sharing108_w;
logic [12:0] sharing109_r, sharing109_w;
logic [12:0] sharing110_r, sharing110_w;
logic [12:0] sharing111_r, sharing111_w;
logic [12:0] sharing112_r, sharing112_w;
logic [12:0] sharing113_r, sharing113_w;
logic [12:0] sharing114_r, sharing114_w;
logic [12:0] sharing115_r, sharing115_w;
logic [12:0] sharing116_r, sharing116_w;
logic [12:0] sharing117_r, sharing117_w;
logic [12:0] sharing118_r, sharing118_w;
logic [12:0] sharing119_r, sharing119_w;
logic [12:0] sharing120_r, sharing120_w;
logic [12:0] sharing121_r, sharing121_w;
logic [12:0] sharing122_r, sharing122_w;
logic [12:0] sharing123_r, sharing123_w;
logic [12:0] sharing124_r, sharing124_w;
logic [12:0] sharing125_r, sharing125_w;
logic [12:0] sharing126_r, sharing126_w;
logic [12:0] sharing127_r, sharing127_w;
logic [12:0] sharing128_r, sharing128_w;
logic [12:0] sharing129_r, sharing129_w;
logic [12:0] sharing130_r, sharing130_w;
logic [12:0] sharing131_r, sharing131_w;
logic [12:0] sharing132_r, sharing132_w;
logic [12:0] sharing133_r, sharing133_w;
logic [12:0] sharing134_r, sharing134_w;
logic [12:0] sharing135_r, sharing135_w;
logic [12:0] sharing136_r, sharing136_w;
logic [12:0] sharing137_r, sharing137_w;
logic [12:0] sharing138_r, sharing138_w;
logic [12:0] sharing139_r, sharing139_w;
logic [12:0] sharing140_r, sharing140_w;
logic [12:0] sharing141_r, sharing141_w;
logic [12:0] sharing142_r, sharing142_w;
logic [12:0] sharing143_r, sharing143_w;
logic [12:0] sharing144_r, sharing144_w;
logic [12:0] sharing145_r, sharing145_w;
logic [12:0] sharing146_r, sharing146_w;
logic [12:0] sharing147_r, sharing147_w;
logic [12:0] sharing148_r, sharing148_w;
logic [12:0] sharing149_r, sharing149_w;
logic [12:0] sharing150_r, sharing150_w;
logic [12:0] sharing151_r, sharing151_w;
logic [12:0] sharing152_r, sharing152_w;
logic [12:0] sharing153_r, sharing153_w;
logic [12:0] sharing154_r, sharing154_w;
logic [12:0] sharing155_r, sharing155_w;
logic [12:0] sharing156_r, sharing156_w;
logic [12:0] sharing157_r, sharing157_w;
logic [12:0] sharing158_r, sharing158_w;
logic [12:0] sharing159_r, sharing159_w;
logic [12:0] sharing160_r, sharing160_w;
logic [12:0] sharing161_r, sharing161_w;
logic [12:0] sharing162_r, sharing162_w;
logic [12:0] sharing163_r, sharing163_w;
logic [12:0] sharing164_r, sharing164_w;
logic [12:0] sharing165_r, sharing165_w;
logic [12:0] sharing166_r, sharing166_w;
logic [12:0] sharing167_r, sharing167_w;
logic [12:0] sharing168_r, sharing168_w;

always_comb begin
	sharing0_w = $signed({in[0],2'b0})+$signed(in[0])+$signed({in[1],2'b0})+$signed(in[57]);
	sharing1_w = $signed({in[2],2'b0})+$signed(in[2])+$signed({in[3],2'b0})+$signed(in[59]);
	sharing2_w = $signed({in[4],2'b0})+$signed(in[4])+$signed({in[5],2'b0})+$signed(in[61]);
	sharing3_w = $signed({in[6],2'b0})+$signed(in[6])+$signed({in[7],2'b0})+$signed(in[63]);
	sharing4_w = $signed({in[8],2'b0})+$signed(in[8])+$signed({in[9],2'b0})+$signed(in[65]);
	sharing5_w = $signed({in[10],2'b0})+$signed(in[10])+$signed({in[11],2'b0})+$signed(in[67]);
	sharing6_w = $signed({in[14],2'b0})+$signed(in[14])+$signed({in[15],2'b0})+$signed(in[71]);
	sharing7_w = $signed({in[16],2'b0})+$signed(in[16])+$signed({in[17],2'b0})+$signed(in[73]);
	sharing8_w = $signed({in[18],2'b0})+$signed(in[18])+$signed({in[19],2'b0})+$signed(in[75]);
	sharing9_w = $signed({in[20],2'b0})+$signed(in[20])+$signed({in[21],2'b0})+$signed(in[77]);
	sharing10_w = $signed({in[22],2'b0})+$signed(in[22])+$signed({in[23],2'b0})+$signed(in[79]);
	sharing11_w = $signed({in[24],2'b0})+$signed(in[24])+$signed({in[25],2'b0})+$signed(in[81]);
	sharing12_w = $signed({in[56],2'b0})+$signed(in[56])+$signed({in[57],2'b0})+$signed(in[113]);
	sharing13_w = $signed({in[60],2'b0})+$signed(in[60])+$signed({in[61],2'b0})+$signed(in[117]);
	sharing14_w = $signed({in[62],2'b0})+$signed(in[62])+$signed({in[63],2'b0})+$signed(in[119]);
	sharing15_w = $signed({in[64],2'b0})+$signed(in[64])+$signed({in[65],2'b0})+$signed(in[121]);
	sharing16_w = $signed({in[66],2'b0})+$signed(in[66])+$signed({in[67],2'b0})+$signed(in[123]);
	sharing17_w = $signed({in[68],2'b0})+$signed(in[68])+$signed({in[69],2'b0})+$signed(in[125]);
	sharing18_w = $signed({in[70],2'b0})+$signed(in[70])+$signed({in[71],2'b0})+$signed(in[127]);
	sharing19_w = $signed({in[72],2'b0})+$signed(in[72])+$signed({in[73],2'b0})+$signed(in[129]);
	sharing20_w = $signed({in[76],2'b0})+$signed(in[76])+$signed({in[77],2'b0})+$signed(in[133]);
	sharing21_w = $signed({in[78],2'b0})+$signed(in[78])+$signed({in[79],2'b0})+$signed(in[135]);
	sharing22_w = $signed({in[80],2'b0})+$signed(in[80])+$signed({in[81],2'b0})+$signed(in[137]);
	sharing23_w = $signed({in[112],2'b0})+$signed(in[112])+$signed({in[113],2'b0})+$signed(in[169]);
	sharing24_w = $signed({in[114],2'b0})+$signed(in[114])+$signed({in[115],2'b0})+$signed(in[171]);
	sharing25_w = $signed({in[116],2'b0})+$signed(in[116])+$signed({in[117],2'b0})+$signed(in[173]);
	sharing26_w = $signed({in[118],2'b0})+$signed(in[118])+$signed({in[119],2'b0})+$signed(in[175]);
	sharing27_w = $signed({in[122],2'b0})+$signed(in[122])+$signed({in[123],2'b0})+$signed(in[179]);
	sharing28_w = $signed({in[124],2'b0})+$signed(in[124])+$signed({in[125],2'b0})+$signed(in[181]);
	sharing29_w = $signed({in[126],2'b0})+$signed(in[126])+$signed({in[127],2'b0})+$signed(in[183]);
	sharing30_w = $signed({in[128],2'b0})+$signed(in[128])+$signed({in[129],2'b0})+$signed(in[185]);
	sharing31_w = $signed({in[130],2'b0})+$signed(in[130])+$signed({in[131],2'b0})+$signed(in[187]);
	sharing32_w = $signed({in[132],2'b0})+$signed(in[132])+$signed({in[133],2'b0})+$signed(in[189]);
	sharing33_w = $signed({in[134],2'b0})+$signed(in[134])+$signed({in[135],2'b0})+$signed(in[191]);
	sharing34_w = $signed({in[168],2'b0})+$signed(in[168])+$signed({in[169],2'b0})+$signed(in[225]);
	sharing35_w = $signed({in[170],2'b0})+$signed(in[170])+$signed({in[171],2'b0})+$signed(in[227]);
	sharing36_w = $signed({in[172],2'b0})+$signed(in[172])+$signed({in[173],2'b0})+$signed(in[229]);
	sharing37_w = $signed({in[174],2'b0})+$signed(in[174])+$signed({in[175],2'b0})+$signed(in[231]);
	sharing38_w = $signed({in[176],2'b0})+$signed(in[176])+$signed({in[177],2'b0})+$signed(in[233]);
	sharing39_w = $signed({in[178],2'b0})+$signed(in[178])+$signed({in[179],2'b0})+$signed(in[235]);
	sharing40_w = $signed({in[180],2'b0})+$signed(in[180])+$signed({in[181],2'b0})+$signed(in[237]);
	sharing41_w = $signed({in[184],2'b0})+$signed(in[184])+$signed({in[185],2'b0})+$signed(in[241]);
	sharing42_w = $signed({in[186],2'b0})+$signed(in[186])+$signed({in[187],2'b0})+$signed(in[243]);
	sharing43_w = $signed({in[188],2'b0})+$signed(in[188])+$signed({in[189],2'b0})+$signed(in[245]);
	sharing44_w = $signed({in[190],2'b0})+$signed(in[190])+$signed({in[191],2'b0})+$signed(in[247]);
	sharing45_w = $signed({in[192],2'b0})+$signed(in[192])+$signed({in[193],2'b0})+$signed(in[249]);
	sharing46_w = $signed({in[224],2'b0})+$signed(in[224])+$signed({in[225],2'b0})+$signed(in[281]);
	sharing47_w = $signed({in[226],2'b0})+$signed(in[226])+$signed({in[227],2'b0})+$signed(in[283]);
	sharing48_w = $signed({in[230],2'b0})+$signed(in[230])+$signed({in[231],2'b0})+$signed(in[287]);
	sharing49_w = $signed({in[232],2'b0})+$signed(in[232])+$signed({in[233],2'b0})+$signed(in[289]);
	sharing50_w = $signed({in[234],2'b0})+$signed(in[234])+$signed({in[235],2'b0})+$signed(in[291]);
	sharing51_w = $signed({in[236],2'b0})+$signed(in[236])+$signed({in[237],2'b0})+$signed(in[293]);
	sharing52_w = $signed({in[238],2'b0})+$signed(in[238])+$signed({in[239],2'b0})+$signed(in[295]);
	sharing53_w = $signed({in[240],2'b0})+$signed(in[240])+$signed({in[241],2'b0})+$signed(in[297]);
	sharing54_w = $signed({in[242],2'b0})+$signed(in[242])+$signed({in[243],2'b0})+$signed(in[299]);
	sharing55_w = $signed({in[246],2'b0})+$signed(in[246])+$signed({in[247],2'b0})+$signed(in[303]);
	sharing56_w = $signed({in[248],2'b0})+$signed(in[248])+$signed({in[249],2'b0})+$signed(in[305]);
	sharing57_w = $signed({in[280],2'b0})+$signed(in[280])+$signed({in[281],2'b0})+$signed(in[337]);
	sharing58_w = $signed({in[282],2'b0})+$signed(in[282])+$signed({in[283],2'b0})+$signed(in[339]);
	sharing59_w = $signed({in[284],2'b0})+$signed(in[284])+$signed({in[285],2'b0})+$signed(in[341]);
	sharing60_w = $signed({in[286],2'b0})+$signed(in[286])+$signed({in[287],2'b0})+$signed(in[343]);
	sharing61_w = $signed({in[288],2'b0})+$signed(in[288])+$signed({in[289],2'b0})+$signed(in[345]);
	sharing62_w = $signed({in[292],2'b0})+$signed(in[292])+$signed({in[293],2'b0})+$signed(in[349]);
	sharing63_w = $signed({in[294],2'b0})+$signed(in[294])+$signed({in[295],2'b0})+$signed(in[351]);
	sharing64_w = $signed({in[296],2'b0})+$signed(in[296])+$signed({in[297],2'b0})+$signed(in[353]);
	sharing65_w = $signed({in[298],2'b0})+$signed(in[298])+$signed({in[299],2'b0})+$signed(in[355]);
	sharing66_w = $signed({in[300],2'b0})+$signed(in[300])+$signed({in[301],2'b0})+$signed(in[357]);
	sharing67_w = $signed({in[302],2'b0})+$signed(in[302])+$signed({in[303],2'b0})+$signed(in[359]);
	sharing68_w = $signed({in[304],2'b0})+$signed(in[304])+$signed({in[305],2'b0})+$signed(in[361]);
	sharing69_w = $signed({in[338],2'b0})+$signed(in[338])+$signed({in[339],2'b0})+$signed(in[395]);
	sharing70_w = $signed({in[340],2'b0})+$signed(in[340])+$signed({in[341],2'b0})+$signed(in[397]);
	sharing71_w = $signed({in[342],2'b0})+$signed(in[342])+$signed({in[343],2'b0})+$signed(in[399]);
	sharing72_w = $signed({in[344],2'b0})+$signed(in[344])+$signed({in[345],2'b0})+$signed(in[401]);
	sharing73_w = $signed({in[346],2'b0})+$signed(in[346])+$signed({in[347],2'b0})+$signed(in[403]);
	sharing74_w = $signed({in[348],2'b0})+$signed(in[348])+$signed({in[349],2'b0})+$signed(in[405]);
	sharing75_w = $signed({in[350],2'b0})+$signed(in[350])+$signed({in[351],2'b0})+$signed(in[407]);
	sharing76_w = $signed({in[354],2'b0})+$signed(in[354])+$signed({in[355],2'b0})+$signed(in[411]);
	sharing77_w = $signed({in[356],2'b0})+$signed(in[356])+$signed({in[357],2'b0})+$signed(in[413]);
	sharing78_w = $signed({in[358],2'b0})+$signed(in[358])+$signed({in[359],2'b0})+$signed(in[415]);
	sharing79_w = $signed({in[360],2'b0})+$signed(in[360])+$signed({in[361],2'b0})+$signed(in[417]);
	sharing80_w = $signed({in[392],2'b0})+$signed(in[392])+$signed({in[393],2'b0})+$signed(in[449]);
	sharing81_w = $signed({in[394],2'b0})+$signed(in[394])+$signed({in[395],2'b0})+$signed(in[451]);
	sharing82_w = $signed({in[396],2'b0})+$signed(in[396])+$signed({in[397],2'b0})+$signed(in[453]);
	sharing83_w = $signed({in[400],2'b0})+$signed(in[400])+$signed({in[401],2'b0})+$signed(in[457]);
	sharing84_w = $signed({in[402],2'b0})+$signed(in[402])+$signed({in[403],2'b0})+$signed(in[459]);
	sharing85_w = $signed({in[404],2'b0})+$signed(in[404])+$signed({in[405],2'b0})+$signed(in[461]);
	sharing86_w = $signed({in[406],2'b0})+$signed(in[406])+$signed({in[407],2'b0})+$signed(in[463]);
	sharing87_w = $signed({in[408],2'b0})+$signed(in[408])+$signed({in[409],2'b0})+$signed(in[465]);
	sharing88_w = $signed({in[410],2'b0})+$signed(in[410])+$signed({in[411],2'b0})+$signed(in[467]);
	sharing89_w = $signed({in[412],2'b0})+$signed(in[412])+$signed({in[413],2'b0})+$signed(in[469]);
	sharing90_w = $signed({in[416],2'b0})+$signed(in[416])+$signed({in[417],2'b0})+$signed(in[473]);
	sharing91_w = $signed({in[448],2'b0})+$signed(in[448])+$signed({in[449],2'b0})+$signed(in[505]);
	sharing92_w = $signed({in[450],2'b0})+$signed(in[450])+$signed({in[451],2'b0})+$signed(in[507]);
	sharing93_w = $signed({in[452],2'b0})+$signed(in[452])+$signed({in[453],2'b0})+$signed(in[509]);
	sharing94_w = $signed({in[454],2'b0})+$signed(in[454])+$signed({in[455],2'b0})+$signed(in[511]);
	sharing95_w = $signed({in[456],2'b0})+$signed(in[456])+$signed({in[457],2'b0})+$signed(in[513]);
	sharing96_w = $signed({in[458],2'b0})+$signed(in[458])+$signed({in[459],2'b0})+$signed(in[515]);
	sharing97_w = $signed({in[462],2'b0})+$signed(in[462])+$signed({in[463],2'b0})+$signed(in[519]);
	sharing98_w = $signed({in[464],2'b0})+$signed(in[464])+$signed({in[465],2'b0})+$signed(in[521]);
	sharing99_w = $signed({in[466],2'b0})+$signed(in[466])+$signed({in[467],2'b0})+$signed(in[523]);
	sharing100_w = $signed({in[468],2'b0})+$signed(in[468])+$signed({in[469],2'b0})+$signed(in[525]);
	sharing101_w = $signed({in[470],2'b0})+$signed(in[470])+$signed({in[471],2'b0})+$signed(in[527]);
	sharing102_w = $signed({in[472],2'b0})+$signed(in[472])+$signed({in[473],2'b0})+$signed(in[529]);
	sharing103_w = $signed({in[504],2'b0})+$signed(in[504])+$signed({in[505],2'b0})+$signed(in[561]);
	sharing104_w = $signed({in[508],2'b0})+$signed(in[508])+$signed({in[509],2'b0})+$signed(in[565]);
	sharing105_w = $signed({in[510],2'b0})+$signed(in[510])+$signed({in[511],2'b0})+$signed(in[567]);
	sharing106_w = $signed({in[512],2'b0})+$signed(in[512])+$signed({in[513],2'b0})+$signed(in[569]);
	sharing107_w = $signed({in[514],2'b0})+$signed(in[514])+$signed({in[515],2'b0})+$signed(in[571]);
	sharing108_w = $signed({in[516],2'b0})+$signed(in[516])+$signed({in[517],2'b0})+$signed(in[573]);
	sharing109_w = $signed({in[518],2'b0})+$signed(in[518])+$signed({in[519],2'b0})+$signed(in[575]);
	sharing110_w = $signed({in[520],2'b0})+$signed(in[520])+$signed({in[521],2'b0})+$signed(in[577]);
	sharing111_w = $signed({in[524],2'b0})+$signed(in[524])+$signed({in[525],2'b0})+$signed(in[581]);
	sharing112_w = $signed({in[526],2'b0})+$signed(in[526])+$signed({in[527],2'b0})+$signed(in[583]);
	sharing113_w = $signed({in[528],2'b0})+$signed(in[528])+$signed({in[529],2'b0})+$signed(in[585]);
	sharing114_w = $signed({in[560],2'b0})+$signed(in[560])+$signed({in[561],2'b0})+$signed(in[617]);
	sharing115_w = $signed({in[562],2'b0})+$signed(in[562])+$signed({in[563],2'b0})+$signed(in[619]);
	sharing116_w = $signed({in[564],2'b0})+$signed(in[564])+$signed({in[565],2'b0})+$signed(in[621]);
	sharing117_w = $signed({in[566],2'b0})+$signed(in[566])+$signed({in[567],2'b0})+$signed(in[623]);
	sharing118_w = $signed({in[570],2'b0})+$signed(in[570])+$signed({in[571],2'b0})+$signed(in[627]);
	sharing119_w = $signed({in[572],2'b0})+$signed(in[572])+$signed({in[573],2'b0})+$signed(in[629]);
	sharing120_w = $signed({in[574],2'b0})+$signed(in[574])+$signed({in[575],2'b0})+$signed(in[631]);
	sharing121_w = $signed({in[576],2'b0})+$signed(in[576])+$signed({in[577],2'b0})+$signed(in[633]);
	sharing122_w = $signed({in[578],2'b0})+$signed(in[578])+$signed({in[579],2'b0})+$signed(in[635]);
	sharing123_w = $signed({in[580],2'b0})+$signed(in[580])+$signed({in[581],2'b0})+$signed(in[637]);
	sharing124_w = $signed({in[582],2'b0})+$signed(in[582])+$signed({in[583],2'b0})+$signed(in[639]);
	sharing125_w = $signed({in[616],2'b0})+$signed(in[616])+$signed({in[617],2'b0})+$signed(in[673]);
	sharing126_w = $signed({in[618],2'b0})+$signed(in[618])+$signed({in[619],2'b0})+$signed(in[675]);
	sharing127_w = $signed({in[620],2'b0})+$signed(in[620])+$signed({in[621],2'b0})+$signed(in[677]);
	sharing128_w = $signed({in[622],2'b0})+$signed(in[622])+$signed({in[623],2'b0})+$signed(in[679]);
	sharing129_w = $signed({in[624],2'b0})+$signed(in[624])+$signed({in[625],2'b0})+$signed(in[681]);
	sharing130_w = $signed({in[626],2'b0})+$signed(in[626])+$signed({in[627],2'b0})+$signed(in[683]);
	sharing131_w = $signed({in[628],2'b0})+$signed(in[628])+$signed({in[629],2'b0})+$signed(in[685]);
	sharing132_w = $signed({in[632],2'b0})+$signed(in[632])+$signed({in[633],2'b0})+$signed(in[689]);
	sharing133_w = $signed({in[634],2'b0})+$signed(in[634])+$signed({in[635],2'b0})+$signed(in[691]);
	sharing134_w = $signed({in[636],2'b0})+$signed(in[636])+$signed({in[637],2'b0})+$signed(in[693]);
	sharing135_w = $signed({in[638],2'b0})+$signed(in[638])+$signed({in[639],2'b0})+$signed(in[695]);
	sharing136_w = $signed({in[640],2'b0})+$signed(in[640])+$signed({in[641],2'b0})+$signed(in[697]);
	sharing137_w = $signed({in[672],2'b0})+$signed(in[672])+$signed({in[673],2'b0})+$signed(in[729]);
	sharing138_w = $signed({in[674],2'b0})+$signed(in[674])+$signed({in[675],2'b0})+$signed(in[731]);
	sharing139_w = $signed({in[678],2'b0})+$signed(in[678])+$signed({in[679],2'b0})+$signed(in[735]);
	sharing140_w = $signed({in[680],2'b0})+$signed(in[680])+$signed({in[681],2'b0})+$signed(in[737]);
	sharing141_w = $signed({in[682],2'b0})+$signed(in[682])+$signed({in[683],2'b0})+$signed(in[739]);
	sharing142_w = $signed({in[684],2'b0})+$signed(in[684])+$signed({in[685],2'b0})+$signed(in[741]);
	sharing143_w = $signed({in[686],2'b0})+$signed(in[686])+$signed({in[687],2'b0})+$signed(in[743]);
	sharing144_w = $signed({in[688],2'b0})+$signed(in[688])+$signed({in[689],2'b0})+$signed(in[745]);
	sharing145_w = $signed({in[690],2'b0})+$signed(in[690])+$signed({in[691],2'b0})+$signed(in[747]);
	sharing146_w = $signed({in[694],2'b0})+$signed(in[694])+$signed({in[695],2'b0})+$signed(in[751]);
	sharing147_w = $signed({in[696],2'b0})+$signed(in[696])+$signed({in[697],2'b0})+$signed(in[753]);
	sharing148_w = $signed({in[12],2'b0})+$signed(in[12])+$signed({in[13],2'b0})+$signed(in[69]);
	sharing149_w = $signed({in[58],2'b0})+$signed(in[58])+$signed({in[59],2'b0})+$signed(in[115]);
	sharing150_w = $signed({in[74],2'b0})+$signed(in[74])+$signed({in[75],2'b0})+$signed(in[131]);
	sharing151_w = $signed({in[120],2'b0})+$signed(in[120])+$signed({in[121],2'b0})+$signed(in[177]);
	sharing152_w = $signed({in[136],2'b0})+$signed(in[136])+$signed({in[137],2'b0})+$signed(in[193]);
	sharing153_w = $signed({in[182],2'b0})+$signed(in[182])+$signed({in[183],2'b0})+$signed(in[239]);
	sharing154_w = $signed({in[228],2'b0})+$signed(in[228])+$signed({in[229],2'b0})+$signed(in[285]);
	sharing155_w = $signed({in[244],2'b0})+$signed(in[244])+$signed({in[245],2'b0})+$signed(in[301]);
	sharing156_w = $signed({in[290],2'b0})+$signed(in[290])+$signed({in[291],2'b0})+$signed(in[347]);
	sharing157_w = $signed({in[336],2'b0})+$signed(in[336])+$signed({in[337],2'b0})+$signed(in[393]);
	sharing158_w = $signed({in[352],2'b0})+$signed(in[352])+$signed({in[353],2'b0})+$signed(in[409]);
	sharing159_w = $signed({in[398],2'b0})+$signed(in[398])+$signed({in[399],2'b0})+$signed(in[455]);
	sharing160_w = $signed({in[414],2'b0})+$signed(in[414])+$signed({in[415],2'b0})+$signed(in[471]);
	sharing161_w = $signed({in[460],2'b0})+$signed(in[460])+$signed({in[461],2'b0})+$signed(in[517]);
	sharing162_w = $signed({in[506],2'b0})+$signed(in[506])+$signed({in[507],2'b0})+$signed(in[563]);
	sharing163_w = $signed({in[522],2'b0})+$signed(in[522])+$signed({in[523],2'b0})+$signed(in[579]);
	sharing164_w = $signed({in[568],2'b0})+$signed(in[568])+$signed({in[569],2'b0})+$signed(in[625]);
	sharing165_w = $signed({in[584],2'b0})+$signed(in[584])+$signed({in[585],2'b0})+$signed(in[641]);
	sharing166_w = $signed({in[630],2'b0})+$signed(in[630])+$signed({in[631],2'b0})+$signed(in[687]);
	sharing167_w = $signed({in[676],2'b0})+$signed(in[676])+$signed({in[677],2'b0})+$signed(in[733]);
	sharing168_w = $signed({in[692],2'b0})+$signed(in[692])+$signed({in[693],2'b0})+$signed(in[749]);
end

assign weighted_sum[0] = $signed(in[0])+$signed(-in[56])+$signed(in[1])+$signed({in[28],2'b0})+$signed(in[28])+$signed({in[29],1'b0})+$signed(in[29])+$signed({in[30],2'b0})+$signed(7);
assign weighted_sum[1] = $signed({in[32],2'b0})+$signed(in[2])+$signed(-in[58])+$signed(in[3])+$signed({in[30],2'b0})+$signed(in[30])+$signed({in[31],1'b0})+$signed(in[31])+$signed(7);
assign weighted_sum[2] = $signed({in[32],2'b0})+$signed(in[32])+$signed({in[33],1'b0})+$signed(in[33])+$signed({in[34],2'b0})+$signed(in[4])+$signed(-in[60])+$signed(in[5])+$signed(7);
assign weighted_sum[3] = $signed(in[6])+$signed({in[34],2'b0})+$signed(in[34])+$signed({in[35],1'b0})+$signed(in[35])+$signed({in[36],2'b0})+$signed(-in[62])+$signed(in[7])+$signed(7);
assign weighted_sum[4] = $signed(-in[64])+$signed(in[8])+$signed(in[9])+$signed({in[36],2'b0})+$signed(in[36])+$signed({in[37],1'b0})+$signed(in[37])+$signed({in[38],2'b0})+$signed(7);
assign weighted_sum[5] = $signed({in[40],2'b0})+$signed(-in[66])+$signed(in[10])+$signed(in[11])+$signed({in[38],2'b0})+$signed(in[38])+$signed({in[39],1'b0})+$signed(in[39])+$signed(7);
assign weighted_sum[6] = $signed({in[40],2'b0})+$signed(in[40])+$signed({in[41],1'b0})+$signed(in[41])+$signed({in[42],2'b0})+$signed(in[12])+$signed(-in[68])+$signed(in[13])+$signed(7);
assign weighted_sum[7] = $signed({in[42],2'b0})+$signed(in[14])+$signed(in[42])+$signed({in[43],1'b0})+$signed(in[43])+$signed({in[44],2'b0})+$signed(-in[70])+$signed(in[15])+$signed(7);
assign weighted_sum[8] = $signed(-in[72])+$signed(in[16])+$signed(in[17])+$signed({in[44],2'b0})+$signed(in[44])+$signed({in[45],1'b0})+$signed(in[45])+$signed({in[46],2'b0})+$signed(7);
assign weighted_sum[9] = $signed({in[48],2'b0})+$signed(in[18])+$signed(-in[74])+$signed(in[19])+$signed({in[46],2'b0})+$signed(in[46])+$signed({in[47],1'b0})+$signed(in[47])+$signed(7);
assign weighted_sum[10] = $signed({in[48],2'b0})+$signed(in[48])+$signed({in[49],1'b0})+$signed(in[49])+$signed({in[50],2'b0})+$signed(in[20])+$signed(-in[76])+$signed(in[21])+$signed(7);
assign weighted_sum[11] = $signed({in[50],2'b0})+$signed(in[22])+$signed(in[50])+$signed({in[51],1'b0})+$signed(in[51])+$signed({in[52],2'b0})+$signed(-in[78])+$signed(in[23])+$signed(7);
assign weighted_sum[12] = $signed(-in[80])+$signed(in[24])+$signed(in[25])+$signed({in[52],2'b0})+$signed(in[52])+$signed({in[53],1'b0})+$signed(in[53])+$signed({in[54],2'b0})+$signed(7);
assign weighted_sum[13] = $signed(in[56])+$signed(-in[112])+$signed(in[57])+$signed({in[84],2'b0})+$signed(in[84])+$signed({in[85],1'b0})+$signed(in[85])+$signed({in[86],2'b0})+$signed(7);
assign weighted_sum[14] = $signed({in[88],2'b0})+$signed(in[58])+$signed(-in[114])+$signed(in[59])+$signed({in[86],2'b0})+$signed(in[86])+$signed({in[87],1'b0})+$signed(in[87])+$signed(7);
assign weighted_sum[15] = $signed({in[88],2'b0})+$signed(in[88])+$signed({in[89],1'b0})+$signed(in[89])+$signed({in[90],2'b0})+$signed(in[60])+$signed(-in[116])+$signed(in[61])+$signed(7);
assign weighted_sum[16] = $signed({in[90],2'b0})+$signed(in[90])+$signed({in[91],1'b0})+$signed(in[91])+$signed(in[62])+$signed({in[92],2'b0})+$signed(-in[118])+$signed(in[63])+$signed(7);
assign weighted_sum[17] = $signed(in[64])+$signed(-in[120])+$signed(in[65])+$signed({in[92],2'b0})+$signed(in[92])+$signed({in[93],1'b0})+$signed(in[93])+$signed({in[94],2'b0})+$signed(7);
assign weighted_sum[18] = $signed({in[96],2'b0})+$signed(in[66])+$signed(-in[122])+$signed(in[67])+$signed({in[94],2'b0})+$signed(in[94])+$signed({in[95],1'b0})+$signed(in[95])+$signed(7);
assign weighted_sum[19] = $signed({in[96],2'b0})+$signed(in[96])+$signed({in[97],1'b0})+$signed(in[97])+$signed({in[98],2'b0})+$signed(in[68])+$signed(-in[124])+$signed(in[69])+$signed(7);
assign weighted_sum[20] = $signed({in[98],2'b0})+$signed(in[98])+$signed({in[99],1'b0})+$signed(in[99])+$signed(in[70])+$signed({in[100],2'b0})+$signed(-in[126])+$signed(in[71])+$signed(7);
assign weighted_sum[21] = $signed(-in[128])+$signed(in[72])+$signed(in[73])+$signed({in[100],2'b0})+$signed(in[100])+$signed({in[101],1'b0})+$signed(in[101])+$signed({in[102],2'b0})+$signed(7);
assign weighted_sum[22] = $signed({in[104],2'b0})+$signed(-in[130])+$signed(in[74])+$signed(in[75])+$signed({in[102],2'b0})+$signed(in[102])+$signed({in[103],1'b0})+$signed(in[103])+$signed(7);
assign weighted_sum[23] = $signed({in[104],2'b0})+$signed(in[104])+$signed({in[105],1'b0})+$signed(in[105])+$signed({in[106],2'b0})+$signed(in[76])+$signed(-in[132])+$signed(in[77])+$signed(7);
assign weighted_sum[24] = $signed({in[106],2'b0})+$signed(in[106])+$signed({in[107],1'b0})+$signed(in[107])+$signed({in[108],2'b0})+$signed(in[78])+$signed(-in[134])+$signed(in[79])+$signed(7);
assign weighted_sum[25] = $signed(-in[136])+$signed(in[80])+$signed(in[81])+$signed({in[108],2'b0})+$signed(in[108])+$signed({in[109],1'b0})+$signed(in[109])+$signed({in[110],2'b0})+$signed(7);
assign weighted_sum[26] = $signed(in[112])+$signed(-in[168])+$signed(in[113])+$signed({in[140],2'b0})+$signed(in[140])+$signed({in[141],1'b0})+$signed(in[141])+$signed({in[142],2'b0})+$signed(7);
assign weighted_sum[27] = $signed({in[144],2'b0})+$signed(in[114])+$signed(-in[170])+$signed(in[115])+$signed({in[142],2'b0})+$signed(in[142])+$signed({in[143],1'b0})+$signed(in[143])+$signed(7);
assign weighted_sum[28] = $signed({in[144],2'b0})+$signed(in[144])+$signed({in[145],1'b0})+$signed(in[145])+$signed({in[146],2'b0})+$signed(in[116])+$signed(-in[172])+$signed(in[117])+$signed(7);
assign weighted_sum[29] = $signed({in[146],2'b0})+$signed(in[146])+$signed({in[147],1'b0})+$signed(in[147])+$signed({in[148],2'b0})+$signed(in[118])+$signed(-in[174])+$signed(in[119])+$signed(7);
assign weighted_sum[30] = $signed(in[120])+$signed(-in[176])+$signed(in[121])+$signed({in[148],2'b0})+$signed(in[148])+$signed({in[149],1'b0})+$signed(in[149])+$signed({in[150],2'b0})+$signed(7);
assign weighted_sum[31] = $signed({in[152],2'b0})+$signed(in[122])+$signed(-in[178])+$signed(in[123])+$signed({in[150],2'b0})+$signed(in[150])+$signed({in[151],1'b0})+$signed(in[151])+$signed(7);
assign weighted_sum[32] = $signed({in[152],2'b0})+$signed(in[152])+$signed({in[153],1'b0})+$signed(in[153])+$signed({in[154],2'b0})+$signed(in[124])+$signed(-in[180])+$signed(in[125])+$signed(7);
assign weighted_sum[33] = $signed({in[154],2'b0})+$signed(in[154])+$signed({in[155],1'b0})+$signed(in[155])+$signed({in[156],2'b0})+$signed(in[126])+$signed(-in[182])+$signed(in[127])+$signed(7);
assign weighted_sum[34] = $signed(in[128])+$signed(-in[184])+$signed(in[129])+$signed({in[156],2'b0})+$signed(in[156])+$signed({in[157],1'b0})+$signed(in[157])+$signed({in[158],2'b0})+$signed(7);
assign weighted_sum[35] = $signed({in[160],2'b0})+$signed(in[130])+$signed(-in[186])+$signed(in[131])+$signed({in[158],2'b0})+$signed(in[158])+$signed({in[159],1'b0})+$signed(in[159])+$signed(7);
assign weighted_sum[36] = $signed({in[160],2'b0})+$signed(in[160])+$signed({in[161],1'b0})+$signed(in[161])+$signed({in[162],2'b0})+$signed(in[132])+$signed(-in[188])+$signed(in[133])+$signed(7);
assign weighted_sum[37] = $signed({in[162],2'b0})+$signed(in[162])+$signed(in[135])+$signed({in[163],1'b0})+$signed(in[163])+$signed({in[164],2'b0})+$signed(in[134])+$signed(-in[190])+$signed(7);
assign weighted_sum[38] = $signed(-in[192])+$signed(in[136])+$signed(in[137])+$signed({in[164],2'b0})+$signed(in[164])+$signed({in[165],1'b0})+$signed(in[165])+$signed({in[166],2'b0})+$signed(7);
assign weighted_sum[39] = $signed(in[168])+$signed(-in[224])+$signed(in[169])+$signed({in[196],2'b0})+$signed(in[196])+$signed({in[197],1'b0})+$signed(in[197])+$signed({in[198],2'b0})+$signed(7);
assign weighted_sum[40] = $signed({in[200],2'b0})+$signed(in[170])+$signed(-in[226])+$signed(in[171])+$signed({in[198],2'b0})+$signed(in[198])+$signed({in[199],1'b0})+$signed(in[199])+$signed(7);
assign weighted_sum[41] = $signed({in[200],2'b0})+$signed(in[200])+$signed({in[201],1'b0})+$signed(in[201])+$signed({in[202],2'b0})+$signed(in[172])+$signed(-in[228])+$signed(in[173])+$signed(7);
assign weighted_sum[42] = $signed({in[202],2'b0})+$signed(in[202])+$signed({in[203],1'b0})+$signed(in[203])+$signed({in[204],2'b0})+$signed(-in[230])+$signed(in[174])+$signed(in[175])+$signed(7);
assign weighted_sum[43] = $signed(in[176])+$signed(-in[232])+$signed(in[177])+$signed({in[204],2'b0})+$signed(in[204])+$signed({in[205],1'b0})+$signed(in[205])+$signed({in[206],2'b0})+$signed(7);
assign weighted_sum[44] = $signed({in[208],2'b0})+$signed(in[178])+$signed(-in[234])+$signed(in[179])+$signed({in[206],2'b0})+$signed(in[206])+$signed({in[207],1'b0})+$signed(in[207])+$signed(7);
assign weighted_sum[45] = $signed({in[208],2'b0})+$signed(in[208])+$signed({in[209],1'b0})+$signed(in[209])+$signed({in[210],2'b0})+$signed(in[180])+$signed(-in[236])+$signed(in[181])+$signed(7);
assign weighted_sum[46] = $signed({in[210],2'b0})+$signed(in[210])+$signed({in[211],1'b0})+$signed(in[211])+$signed({in[212],2'b0})+$signed(-in[238])+$signed(in[182])+$signed(in[183])+$signed(7);
assign weighted_sum[47] = $signed(in[184])+$signed(-in[240])+$signed(in[185])+$signed({in[212],2'b0})+$signed(in[212])+$signed({in[213],1'b0})+$signed(in[213])+$signed({in[214],2'b0})+$signed(7);
assign weighted_sum[48] = $signed({in[216],2'b0})+$signed(in[186])+$signed(-in[242])+$signed(in[187])+$signed({in[214],2'b0})+$signed(in[214])+$signed({in[215],1'b0})+$signed(in[215])+$signed(7);
assign weighted_sum[49] = $signed({in[216],2'b0})+$signed(in[216])+$signed({in[217],1'b0})+$signed(in[217])+$signed({in[218],2'b0})+$signed(in[188])+$signed(-in[244])+$signed(in[189])+$signed(7);
assign weighted_sum[50] = $signed({in[218],2'b0})+$signed(in[218])+$signed({in[219],1'b0})+$signed(in[219])+$signed({in[220],2'b0})+$signed(in[191])+$signed(-in[246])+$signed(in[190])+$signed(7);
assign weighted_sum[51] = $signed(in[192])+$signed(-in[248])+$signed(in[193])+$signed({in[220],2'b0})+$signed(in[220])+$signed({in[221],1'b0})+$signed(in[221])+$signed({in[222],2'b0})+$signed(7);
assign weighted_sum[52] = $signed(-in[280])+$signed(in[224])+$signed(in[225])+$signed({in[252],2'b0})+$signed(in[252])+$signed({in[253],1'b0})+$signed(in[253])+$signed({in[254],2'b0})+$signed(7);
assign weighted_sum[53] = $signed({in[256],2'b0})+$signed(in[226])+$signed(-in[282])+$signed(in[227])+$signed({in[254],2'b0})+$signed(in[254])+$signed({in[255],1'b0})+$signed(in[255])+$signed(7);
assign weighted_sum[54] = $signed({in[256],2'b0})+$signed(in[256])+$signed({in[257],1'b0})+$signed(in[257])+$signed({in[258],2'b0})+$signed(in[228])+$signed(-in[284])+$signed(in[229])+$signed(7);
assign weighted_sum[55] = $signed(in[230])+$signed({in[258],2'b0})+$signed(in[258])+$signed({in[259],1'b0})+$signed(in[259])+$signed({in[260],2'b0})+$signed(-in[286])+$signed(in[231])+$signed(7);
assign weighted_sum[56] = $signed(in[232])+$signed(-in[288])+$signed(in[233])+$signed({in[260],2'b0})+$signed(in[260])+$signed({in[261],1'b0})+$signed(in[261])+$signed({in[262],2'b0})+$signed(7);
assign weighted_sum[57] = $signed({in[264],2'b0})+$signed(in[234])+$signed(-in[290])+$signed(in[235])+$signed({in[262],2'b0})+$signed(in[262])+$signed({in[263],1'b0})+$signed(in[263])+$signed(7);
assign weighted_sum[58] = $signed({in[264],2'b0})+$signed(in[264])+$signed({in[265],1'b0})+$signed(in[265])+$signed({in[266],2'b0})+$signed(in[236])+$signed(-in[292])+$signed(in[237])+$signed(7);
assign weighted_sum[59] = $signed(in[238])+$signed({in[266],2'b0})+$signed(in[266])+$signed({in[267],1'b0})+$signed(in[267])+$signed({in[268],2'b0})+$signed(-in[294])+$signed(in[239])+$signed(7);
assign weighted_sum[60] = $signed(in[240])+$signed(-in[296])+$signed(in[241])+$signed({in[268],2'b0})+$signed(in[268])+$signed({in[269],1'b0})+$signed(in[269])+$signed({in[270],2'b0})+$signed(7);
assign weighted_sum[61] = $signed({in[272],2'b0})+$signed(in[242])+$signed(-in[298])+$signed(in[243])+$signed({in[270],2'b0})+$signed(in[270])+$signed({in[271],1'b0})+$signed(in[271])+$signed(7);
assign weighted_sum[62] = $signed({in[272],2'b0})+$signed(in[272])+$signed({in[273],1'b0})+$signed(in[273])+$signed({in[274],2'b0})+$signed(in[244])+$signed(-in[300])+$signed(in[245])+$signed(7);
assign weighted_sum[63] = $signed(in[246])+$signed({in[274],2'b0})+$signed(in[274])+$signed({in[275],1'b0})+$signed(in[275])+$signed({in[276],2'b0})+$signed(-in[302])+$signed(in[247])+$signed(7);
assign weighted_sum[64] = $signed(in[248])+$signed(-in[304])+$signed(in[249])+$signed({in[276],2'b0})+$signed(in[276])+$signed({in[277],1'b0})+$signed(in[277])+$signed({in[278],2'b0})+$signed(7);
assign weighted_sum[65] = $signed(-in[336])+$signed(in[280])+$signed(in[281])+$signed({in[308],2'b0})+$signed(in[308])+$signed({in[309],1'b0})+$signed(in[309])+$signed({in[310],2'b0})+$signed(7);
assign weighted_sum[66] = $signed({in[312],2'b0})+$signed(-in[338])+$signed(in[282])+$signed(in[283])+$signed({in[310],2'b0})+$signed(in[310])+$signed({in[311],1'b0})+$signed(in[311])+$signed(7);
assign weighted_sum[67] = $signed({in[312],2'b0})+$signed(in[312])+$signed({in[313],1'b0})+$signed(in[313])+$signed({in[314],2'b0})+$signed(in[284])+$signed(-in[340])+$signed(in[285])+$signed(7);
assign weighted_sum[68] = $signed({in[314],2'b0})+$signed(in[314])+$signed(in[286])+$signed({in[315],1'b0})+$signed(in[315])+$signed({in[316],2'b0})+$signed(-in[342])+$signed(in[287])+$signed(7);
assign weighted_sum[69] = $signed(-in[344])+$signed(in[288])+$signed(in[289])+$signed({in[316],2'b0})+$signed(in[316])+$signed({in[317],1'b0})+$signed(in[317])+$signed({in[318],2'b0})+$signed(7);
assign weighted_sum[70] = $signed({in[320],2'b0})+$signed(in[290])+$signed(-in[346])+$signed(in[291])+$signed({in[318],2'b0})+$signed(in[318])+$signed({in[319],1'b0})+$signed(in[319])+$signed(7);
assign weighted_sum[71] = $signed({in[320],2'b0})+$signed(in[320])+$signed({in[321],1'b0})+$signed(in[321])+$signed({in[322],2'b0})+$signed(in[292])+$signed(-in[348])+$signed(in[293])+$signed(7);
assign weighted_sum[72] = $signed({in[322],2'b0})+$signed(in[322])+$signed(in[294])+$signed({in[323],1'b0})+$signed(in[323])+$signed({in[324],2'b0})+$signed(-in[350])+$signed(in[295])+$signed(7);
assign weighted_sum[73] = $signed(in[296])+$signed(-in[352])+$signed(in[297])+$signed({in[324],2'b0})+$signed(in[324])+$signed({in[325],1'b0})+$signed(in[325])+$signed({in[326],2'b0})+$signed(7);
assign weighted_sum[74] = $signed({in[328],2'b0})+$signed(in[298])+$signed(-in[354])+$signed(in[299])+$signed({in[326],2'b0})+$signed(in[326])+$signed({in[327],1'b0})+$signed(in[327])+$signed(7);
assign weighted_sum[75] = $signed({in[328],2'b0})+$signed(in[328])+$signed({in[329],1'b0})+$signed(in[329])+$signed({in[330],2'b0})+$signed(in[300])+$signed(-in[356])+$signed(in[301])+$signed(7);
assign weighted_sum[76] = $signed({in[330],2'b0})+$signed(in[330])+$signed(in[302])+$signed({in[331],1'b0})+$signed(in[331])+$signed({in[332],2'b0})+$signed(-in[358])+$signed(in[303])+$signed(7);
assign weighted_sum[77] = $signed(in[304])+$signed(-in[360])+$signed(in[305])+$signed({in[332],2'b0})+$signed(in[332])+$signed({in[333],1'b0})+$signed(in[333])+$signed({in[334],2'b0})+$signed(7);
assign weighted_sum[78] = $signed(-in[392])+$signed(in[336])+$signed(in[337])+$signed({in[364],2'b0})+$signed(in[364])+$signed({in[365],1'b0})+$signed(in[365])+$signed({in[366],2'b0})+$signed(7);
assign weighted_sum[79] = $signed({in[368],2'b0})+$signed(in[338])+$signed(-in[394])+$signed(in[339])+$signed({in[366],2'b0})+$signed(in[366])+$signed({in[367],1'b0})+$signed(in[367])+$signed(7);
assign weighted_sum[80] = $signed({in[368],2'b0})+$signed(in[368])+$signed({in[369],1'b0})+$signed(in[369])+$signed({in[370],2'b0})+$signed(in[340])+$signed(-in[396])+$signed(in[341])+$signed(7);
assign weighted_sum[81] = $signed({in[370],2'b0})+$signed(in[370])+$signed({in[371],1'b0})+$signed(in[371])+$signed({in[372],2'b0})+$signed(in[342])+$signed(-in[398])+$signed(in[343])+$signed(7);
assign weighted_sum[82] = $signed(-in[400])+$signed(in[344])+$signed(in[345])+$signed({in[372],2'b0})+$signed(in[372])+$signed({in[373],1'b0})+$signed(in[373])+$signed({in[374],2'b0})+$signed(7);
assign weighted_sum[83] = $signed({in[376],2'b0})+$signed(-in[402])+$signed(in[346])+$signed(in[347])+$signed({in[374],2'b0})+$signed(in[374])+$signed({in[375],1'b0})+$signed(in[375])+$signed(7);
assign weighted_sum[84] = $signed({in[376],2'b0})+$signed(in[376])+$signed({in[377],1'b0})+$signed(in[377])+$signed({in[378],2'b0})+$signed(in[348])+$signed(-in[404])+$signed(in[349])+$signed(7);
assign weighted_sum[85] = $signed({in[378],2'b0})+$signed(in[378])+$signed({in[379],1'b0})+$signed(in[379])+$signed({in[380],2'b0})+$signed(in[350])+$signed(-in[406])+$signed(in[351])+$signed(7);
assign weighted_sum[86] = $signed(-in[408])+$signed(in[352])+$signed(in[353])+$signed({in[380],2'b0})+$signed(in[380])+$signed({in[381],1'b0})+$signed(in[381])+$signed({in[382],2'b0})+$signed(7);
assign weighted_sum[87] = $signed({in[384],2'b0})+$signed(in[354])+$signed(-in[410])+$signed(in[355])+$signed({in[382],2'b0})+$signed(in[382])+$signed({in[383],1'b0})+$signed(in[383])+$signed(7);
assign weighted_sum[88] = $signed({in[384],2'b0})+$signed(in[384])+$signed({in[385],1'b0})+$signed(in[385])+$signed({in[386],2'b0})+$signed(in[356])+$signed(-in[412])+$signed(in[357])+$signed(7);
assign weighted_sum[89] = $signed({in[386],2'b0})+$signed(in[386])+$signed({in[387],1'b0})+$signed(in[387])+$signed({in[388],2'b0})+$signed(in[358])+$signed(-in[414])+$signed(in[359])+$signed(7);
assign weighted_sum[90] = $signed(in[360])+$signed(-in[416])+$signed(in[361])+$signed({in[388],2'b0})+$signed(in[388])+$signed({in[389],1'b0})+$signed(in[389])+$signed({in[390],2'b0})+$signed(7);
assign weighted_sum[91] = $signed(-in[448])+$signed(in[392])+$signed(in[393])+$signed({in[420],2'b0})+$signed(in[420])+$signed({in[421],1'b0})+$signed(in[421])+$signed({in[422],2'b0})+$signed(7);
assign weighted_sum[92] = $signed({in[424],2'b0})+$signed(-in[450])+$signed(in[394])+$signed(in[395])+$signed({in[422],2'b0})+$signed(in[422])+$signed({in[423],1'b0})+$signed(in[423])+$signed(7);
assign weighted_sum[93] = $signed({in[424],2'b0})+$signed(in[424])+$signed({in[425],1'b0})+$signed(in[425])+$signed({in[426],2'b0})+$signed(in[396])+$signed(-in[452])+$signed(in[397])+$signed(7);
assign weighted_sum[94] = $signed({in[426],2'b0})+$signed(in[426])+$signed({in[427],1'b0})+$signed(in[427])+$signed({in[428],2'b0})+$signed(in[398])+$signed(-in[454])+$signed(in[399])+$signed(7);
assign weighted_sum[95] = $signed(-in[456])+$signed(in[400])+$signed(in[401])+$signed({in[428],2'b0})+$signed(in[428])+$signed({in[429],1'b0})+$signed(in[429])+$signed({in[430],2'b0})+$signed(7);
assign weighted_sum[96] = $signed({in[432],2'b0})+$signed(in[402])+$signed(-in[458])+$signed(in[403])+$signed({in[430],2'b0})+$signed(in[430])+$signed({in[431],1'b0})+$signed(in[431])+$signed(7);
assign weighted_sum[97] = $signed({in[432],2'b0})+$signed(in[432])+$signed({in[433],1'b0})+$signed(in[433])+$signed({in[434],2'b0})+$signed(in[404])+$signed(-in[460])+$signed(in[405])+$signed(7);
assign weighted_sum[98] = $signed({in[434],2'b0})+$signed(in[434])+$signed({in[435],1'b0})+$signed(in[435])+$signed({in[436],2'b0})+$signed(in[406])+$signed(-in[462])+$signed(in[407])+$signed(7);
assign weighted_sum[99] = $signed(-in[464])+$signed(in[408])+$signed(in[409])+$signed({in[436],2'b0})+$signed(in[436])+$signed({in[437],1'b0})+$signed(in[437])+$signed({in[438],2'b0})+$signed(7);
assign weighted_sum[100] = $signed({in[440],2'b0})+$signed(-in[466])+$signed(in[410])+$signed(in[411])+$signed({in[438],2'b0})+$signed(in[438])+$signed({in[439],1'b0})+$signed(in[439])+$signed(7);
assign weighted_sum[101] = $signed({in[440],2'b0})+$signed(in[440])+$signed({in[441],1'b0})+$signed(in[441])+$signed({in[442],2'b0})+$signed(in[412])+$signed(-in[468])+$signed(in[413])+$signed(7);
assign weighted_sum[102] = $signed({in[442],2'b0})+$signed(in[414])+$signed(in[442])+$signed({in[443],1'b0})+$signed(in[443])+$signed({in[444],2'b0})+$signed(-in[470])+$signed(in[415])+$signed(7);
assign weighted_sum[103] = $signed(-in[472])+$signed(in[416])+$signed(in[417])+$signed({in[444],2'b0})+$signed(in[444])+$signed({in[445],1'b0})+$signed(in[445])+$signed({in[446],2'b0})+$signed(7);
assign weighted_sum[104] = $signed(in[448])+$signed(-in[504])+$signed(in[449])+$signed({in[476],2'b0})+$signed(in[476])+$signed({in[477],1'b0})+$signed(in[477])+$signed({in[478],2'b0})+$signed(7);
assign weighted_sum[105] = $signed({in[480],2'b0})+$signed(in[450])+$signed(-in[506])+$signed(in[451])+$signed({in[478],2'b0})+$signed(in[478])+$signed({in[479],1'b0})+$signed(in[479])+$signed(7);
assign weighted_sum[106] = $signed({in[480],2'b0})+$signed(in[480])+$signed({in[481],1'b0})+$signed(in[481])+$signed({in[482],2'b0})+$signed(in[452])+$signed(-in[508])+$signed(in[453])+$signed(7);
assign weighted_sum[107] = $signed(in[454])+$signed({in[482],2'b0})+$signed(in[482])+$signed({in[483],1'b0})+$signed(in[483])+$signed({in[484],2'b0})+$signed(-in[510])+$signed(in[455])+$signed(7);
assign weighted_sum[108] = $signed(-in[512])+$signed(in[456])+$signed(in[457])+$signed({in[484],2'b0})+$signed(in[484])+$signed({in[485],1'b0})+$signed(in[485])+$signed({in[486],2'b0})+$signed(7);
assign weighted_sum[109] = $signed({in[488],2'b0})+$signed(-in[514])+$signed(in[458])+$signed(in[459])+$signed({in[486],2'b0})+$signed(in[486])+$signed({in[487],1'b0})+$signed(in[487])+$signed(7);
assign weighted_sum[110] = $signed({in[488],2'b0})+$signed(in[488])+$signed({in[489],1'b0})+$signed(in[489])+$signed({in[490],2'b0})+$signed(in[460])+$signed(-in[516])+$signed(in[461])+$signed(7);
assign weighted_sum[111] = $signed(in[462])+$signed({in[490],2'b0})+$signed(in[490])+$signed({in[491],1'b0})+$signed(in[491])+$signed({in[492],2'b0})+$signed(-in[518])+$signed(in[463])+$signed(7);
assign weighted_sum[112] = $signed(-in[520])+$signed(in[464])+$signed(in[465])+$signed({in[492],2'b0})+$signed(in[492])+$signed({in[493],1'b0})+$signed(in[493])+$signed({in[494],2'b0})+$signed(7);
assign weighted_sum[113] = $signed({in[496],2'b0})+$signed(-in[522])+$signed(in[466])+$signed(in[467])+$signed({in[494],2'b0})+$signed(in[494])+$signed({in[495],1'b0})+$signed(in[495])+$signed(7);
assign weighted_sum[114] = $signed({in[496],2'b0})+$signed(in[496])+$signed({in[497],1'b0})+$signed(in[497])+$signed({in[498],2'b0})+$signed(in[468])+$signed(-in[524])+$signed(in[469])+$signed(7);
assign weighted_sum[115] = $signed(in[470])+$signed({in[498],2'b0})+$signed(in[498])+$signed({in[499],1'b0})+$signed(in[499])+$signed({in[500],2'b0})+$signed(-in[526])+$signed(in[471])+$signed(7);
assign weighted_sum[116] = $signed(-in[528])+$signed(in[472])+$signed(in[473])+$signed({in[500],2'b0})+$signed(in[500])+$signed({in[501],1'b0})+$signed(in[501])+$signed({in[502],2'b0})+$signed(7);
assign weighted_sum[117] = $signed(in[504])+$signed(-in[560])+$signed(in[505])+$signed({in[532],2'b0})+$signed(in[532])+$signed({in[533],1'b0})+$signed(in[533])+$signed({in[534],2'b0})+$signed(7);
assign weighted_sum[118] = $signed({in[536],2'b0})+$signed(in[506])+$signed(-in[562])+$signed(in[507])+$signed({in[534],2'b0})+$signed(in[534])+$signed({in[535],1'b0})+$signed(in[535])+$signed(7);
assign weighted_sum[119] = $signed({in[536],2'b0})+$signed(in[536])+$signed({in[537],1'b0})+$signed(in[537])+$signed({in[538],2'b0})+$signed(in[508])+$signed(-in[564])+$signed(in[509])+$signed(7);
assign weighted_sum[120] = $signed(in[510])+$signed({in[538],2'b0})+$signed(in[538])+$signed({in[539],1'b0})+$signed(in[539])+$signed({in[540],2'b0})+$signed(-in[566])+$signed(in[511])+$signed(7);
assign weighted_sum[121] = $signed(in[512])+$signed(-in[568])+$signed(in[513])+$signed({in[540],2'b0})+$signed(in[540])+$signed({in[541],1'b0})+$signed(in[541])+$signed({in[542],2'b0})+$signed(7);
assign weighted_sum[122] = $signed({in[544],2'b0})+$signed(in[514])+$signed(-in[570])+$signed(in[515])+$signed({in[542],2'b0})+$signed(in[542])+$signed({in[543],1'b0})+$signed(in[543])+$signed(7);
assign weighted_sum[123] = $signed({in[544],2'b0})+$signed(in[544])+$signed({in[545],1'b0})+$signed(in[545])+$signed({in[546],2'b0})+$signed(in[516])+$signed(-in[572])+$signed(in[517])+$signed(7);
assign weighted_sum[124] = $signed(in[518])+$signed({in[546],2'b0})+$signed(in[546])+$signed({in[547],1'b0})+$signed(in[547])+$signed({in[548],2'b0})+$signed(-in[574])+$signed(in[519])+$signed(7);
assign weighted_sum[125] = $signed(-in[576])+$signed(in[520])+$signed(in[521])+$signed({in[548],2'b0})+$signed(in[548])+$signed({in[549],1'b0})+$signed(in[549])+$signed({in[550],2'b0})+$signed(7);
assign weighted_sum[126] = $signed({in[552],2'b0})+$signed(-in[578])+$signed(in[522])+$signed(in[523])+$signed({in[550],2'b0})+$signed(in[550])+$signed({in[551],1'b0})+$signed(in[551])+$signed(7);
assign weighted_sum[127] = $signed({in[552],2'b0})+$signed(in[552])+$signed({in[553],1'b0})+$signed(in[553])+$signed({in[554],2'b0})+$signed(in[524])+$signed(-in[580])+$signed(in[525])+$signed(7);
assign weighted_sum[128] = $signed({in[554],2'b0})+$signed(in[526])+$signed(in[554])+$signed({in[555],1'b0})+$signed(in[555])+$signed({in[556],2'b0})+$signed(-in[582])+$signed(in[527])+$signed(7);
assign weighted_sum[129] = $signed(-in[584])+$signed(in[528])+$signed(in[529])+$signed({in[556],2'b0})+$signed(in[556])+$signed({in[557],1'b0})+$signed(in[557])+$signed({in[558],2'b0})+$signed(7);
assign weighted_sum[130] = $signed(in[560])+$signed(-in[616])+$signed(in[561])+$signed({in[588],2'b0})+$signed(in[588])+$signed({in[589],1'b0})+$signed(in[589])+$signed({in[590],2'b0})+$signed(7);
assign weighted_sum[131] = $signed({in[592],2'b0})+$signed(in[562])+$signed(-in[618])+$signed(in[563])+$signed({in[590],2'b0})+$signed(in[590])+$signed({in[591],1'b0})+$signed(in[591])+$signed(7);
assign weighted_sum[132] = $signed({in[592],2'b0})+$signed(in[592])+$signed({in[593],1'b0})+$signed(in[593])+$signed({in[594],2'b0})+$signed(in[564])+$signed(-in[620])+$signed(in[565])+$signed(7);
assign weighted_sum[133] = $signed({in[594],2'b0})+$signed(in[594])+$signed({in[595],1'b0})+$signed(in[595])+$signed(in[566])+$signed({in[596],2'b0})+$signed(-in[622])+$signed(in[567])+$signed(7);
assign weighted_sum[134] = $signed(in[568])+$signed(-in[624])+$signed(in[569])+$signed({in[596],2'b0})+$signed(in[596])+$signed({in[597],1'b0})+$signed(in[597])+$signed({in[598],2'b0})+$signed(7);
assign weighted_sum[135] = $signed({in[600],2'b0})+$signed(in[570])+$signed(-in[626])+$signed(in[571])+$signed({in[598],2'b0})+$signed(in[598])+$signed({in[599],1'b0})+$signed(in[599])+$signed(7);
assign weighted_sum[136] = $signed({in[600],2'b0})+$signed(in[600])+$signed({in[601],1'b0})+$signed(in[601])+$signed({in[602],2'b0})+$signed(in[572])+$signed(-in[628])+$signed(in[573])+$signed(7);
assign weighted_sum[137] = $signed({in[602],2'b0})+$signed(in[602])+$signed({in[603],1'b0})+$signed(in[603])+$signed(in[574])+$signed({in[604],2'b0})+$signed(-in[630])+$signed(in[575])+$signed(7);
assign weighted_sum[138] = $signed(in[576])+$signed(-in[632])+$signed(in[577])+$signed({in[604],2'b0})+$signed(in[604])+$signed({in[605],1'b0})+$signed(in[605])+$signed({in[606],2'b0})+$signed(7);
assign weighted_sum[139] = $signed({in[608],2'b0})+$signed(in[578])+$signed(-in[634])+$signed(in[579])+$signed({in[606],2'b0})+$signed(in[606])+$signed({in[607],1'b0})+$signed(in[607])+$signed(7);
assign weighted_sum[140] = $signed({in[608],2'b0})+$signed(in[608])+$signed({in[609],1'b0})+$signed(in[609])+$signed({in[610],2'b0})+$signed(in[580])+$signed(-in[636])+$signed(in[581])+$signed(7);
assign weighted_sum[141] = $signed({in[610],2'b0})+$signed(in[610])+$signed({in[611],1'b0})+$signed(in[611])+$signed(in[582])+$signed({in[612],2'b0})+$signed(-in[638])+$signed(in[583])+$signed(7);
assign weighted_sum[142] = $signed(-in[640])+$signed(in[584])+$signed(in[585])+$signed({in[612],2'b0})+$signed(in[612])+$signed({in[613],1'b0})+$signed(in[613])+$signed({in[614],2'b0})+$signed(7);
assign weighted_sum[143] = $signed(in[616])+$signed(-in[672])+$signed(in[617])+$signed({in[644],2'b0})+$signed(in[644])+$signed({in[645],1'b0})+$signed(in[645])+$signed({in[646],2'b0})+$signed(7);
assign weighted_sum[144] = $signed({in[648],2'b0})+$signed(in[618])+$signed(-in[674])+$signed(in[619])+$signed({in[646],2'b0})+$signed(in[646])+$signed({in[647],1'b0})+$signed(in[647])+$signed(7);
assign weighted_sum[145] = $signed({in[648],2'b0})+$signed(in[648])+$signed({in[649],1'b0})+$signed(in[649])+$signed({in[650],2'b0})+$signed(in[620])+$signed(-in[676])+$signed(in[621])+$signed(7);
assign weighted_sum[146] = $signed({in[650],2'b0})+$signed(in[650])+$signed({in[651],1'b0})+$signed(in[651])+$signed({in[652],2'b0})+$signed(in[622])+$signed(-in[678])+$signed(in[623])+$signed(7);
assign weighted_sum[147] = $signed(in[624])+$signed(-in[680])+$signed(in[625])+$signed({in[652],2'b0})+$signed(in[652])+$signed({in[653],1'b0})+$signed(in[653])+$signed({in[654],2'b0})+$signed(7);
assign weighted_sum[148] = $signed({in[656],2'b0})+$signed(in[626])+$signed(-in[682])+$signed(in[627])+$signed({in[654],2'b0})+$signed(in[654])+$signed({in[655],1'b0})+$signed(in[655])+$signed(7);
assign weighted_sum[149] = $signed({in[656],2'b0})+$signed(in[656])+$signed({in[657],1'b0})+$signed(in[657])+$signed({in[658],2'b0})+$signed(in[628])+$signed(-in[684])+$signed(in[629])+$signed(7);
assign weighted_sum[150] = $signed({in[658],2'b0})+$signed(in[658])+$signed({in[659],1'b0})+$signed(in[659])+$signed({in[660],2'b0})+$signed(in[630])+$signed(-in[686])+$signed(in[631])+$signed(7);
assign weighted_sum[151] = $signed(in[632])+$signed(-in[688])+$signed(in[633])+$signed({in[660],2'b0})+$signed(in[660])+$signed({in[661],1'b0})+$signed(in[661])+$signed({in[662],2'b0})+$signed(7);
assign weighted_sum[152] = $signed({in[664],2'b0})+$signed(in[634])+$signed(-in[690])+$signed(in[635])+$signed({in[662],2'b0})+$signed(in[662])+$signed({in[663],1'b0})+$signed(in[663])+$signed(7);
assign weighted_sum[153] = $signed({in[664],2'b0})+$signed(in[664])+$signed({in[665],1'b0})+$signed(in[665])+$signed({in[666],2'b0})+$signed(in[636])+$signed(-in[692])+$signed(in[637])+$signed(7);
assign weighted_sum[154] = $signed({in[666],2'b0})+$signed(in[666])+$signed({in[667],1'b0})+$signed(in[667])+$signed({in[668],2'b0})+$signed(in[638])+$signed(-in[694])+$signed(in[639])+$signed(7);
assign weighted_sum[155] = $signed(in[640])+$signed(-in[696])+$signed(in[641])+$signed({in[668],2'b0})+$signed(in[668])+$signed({in[669],1'b0})+$signed(in[669])+$signed({in[670],2'b0})+$signed(7);
assign weighted_sum[156] = $signed(-in[728])+$signed(in[672])+$signed(in[673])+$signed({in[700],2'b0})+$signed(in[700])+$signed({in[701],1'b0})+$signed(in[701])+$signed({in[702],2'b0})+$signed(7);
assign weighted_sum[157] = $signed({in[704],2'b0})+$signed(-in[730])+$signed(in[674])+$signed(in[675])+$signed({in[702],2'b0})+$signed(in[702])+$signed({in[703],1'b0})+$signed(in[703])+$signed(7);
assign weighted_sum[158] = $signed({in[704],2'b0})+$signed(in[704])+$signed({in[705],1'b0})+$signed(in[705])+$signed({in[706],2'b0})+$signed(in[676])+$signed(-in[732])+$signed(in[677])+$signed(7);
assign weighted_sum[159] = $signed({in[706],2'b0})+$signed(in[706])+$signed({in[707],1'b0})+$signed(in[707])+$signed({in[708],2'b0})+$signed(-in[734])+$signed(in[678])+$signed(in[679])+$signed(7);
assign weighted_sum[160] = $signed(in[680])+$signed(-in[736])+$signed(in[681])+$signed({in[708],2'b0})+$signed(in[708])+$signed({in[709],1'b0})+$signed(in[709])+$signed({in[710],2'b0})+$signed(7);
assign weighted_sum[161] = $signed({in[712],2'b0})+$signed(in[682])+$signed(-in[738])+$signed(in[683])+$signed({in[710],2'b0})+$signed(in[710])+$signed({in[711],1'b0})+$signed(in[711])+$signed(7);
assign weighted_sum[162] = $signed({in[712],2'b0})+$signed(in[712])+$signed({in[713],1'b0})+$signed(in[713])+$signed({in[714],2'b0})+$signed(in[684])+$signed(-in[740])+$signed(in[685])+$signed(7);
assign weighted_sum[163] = $signed({in[714],2'b0})+$signed(in[714])+$signed({in[715],1'b0})+$signed(in[715])+$signed({in[716],2'b0})+$signed(-in[742])+$signed(in[686])+$signed(in[687])+$signed(7);
assign weighted_sum[164] = $signed(in[688])+$signed(-in[744])+$signed(in[689])+$signed({in[716],2'b0})+$signed(in[716])+$signed({in[717],1'b0})+$signed(in[717])+$signed({in[718],2'b0})+$signed(7);
assign weighted_sum[165] = $signed({in[720],2'b0})+$signed(in[690])+$signed(-in[746])+$signed(in[691])+$signed({in[718],2'b0})+$signed(in[718])+$signed({in[719],1'b0})+$signed(in[719])+$signed(7);
assign weighted_sum[166] = $signed({in[720],2'b0})+$signed(in[720])+$signed({in[721],1'b0})+$signed(in[721])+$signed({in[722],2'b0})+$signed(in[692])+$signed(-in[748])+$signed(in[693])+$signed(7);
assign weighted_sum[167] = $signed({in[722],2'b0})+$signed(in[722])+$signed({in[723],1'b0})+$signed(in[723])+$signed({in[724],2'b0})+$signed(-in[750])+$signed(in[694])+$signed(in[695])+$signed(7);
assign weighted_sum[168] = $signed(in[696])+$signed(-in[752])+$signed(in[697])+$signed({in[724],2'b0})+$signed(in[724])+$signed({in[725],1'b0})+$signed(in[725])+$signed({in[726],2'b0})+$signed(7);
assign weighted_sum[169] = $signed({in[56],1'b0})+$signed(-{in[57],2'b0})+$signed(-{in[58],2'b0})+$signed(-in[2])+$signed({in[28],1'b0})+$signed(in[28])+$signed(-{in[30],2'b0})+$signed(sharing0_r)+$signed(1);
assign weighted_sum[170] = $signed(-{in[32],2'b0})+$signed({in[58],1'b0})+$signed(-{in[59],2'b0})+$signed(-{in[60],2'b0})+$signed(-in[4])+$signed({in[30],1'b0})+$signed(in[30])+$signed(sharing1_r)+$signed(1);
assign weighted_sum[171] = $signed({in[32],1'b0})+$signed(in[32])+$signed(-{in[34],2'b0})+$signed({in[60],1'b0})+$signed(-{in[61],2'b0})+$signed(-{in[62],2'b0})+$signed(-in[6])+$signed(sharing2_r)+$signed(1);
assign weighted_sum[172] = $signed(-{in[64],2'b0})+$signed(-in[8])+$signed({in[34],1'b0})+$signed(in[34])+$signed(-{in[36],2'b0})+$signed({in[62],1'b0})+$signed(-{in[63],2'b0})+$signed(sharing3_r)+$signed(1);
assign weighted_sum[173] = $signed({in[64],1'b0})+$signed(-{in[65],2'b0})+$signed(-{in[66],2'b0})+$signed(-in[10])+$signed({in[36],1'b0})+$signed(in[36])+$signed(-{in[38],2'b0})+$signed(sharing4_r)+$signed(1);
assign weighted_sum[174] = $signed(-{in[40],2'b0})+$signed({in[66],1'b0})+$signed(-{in[67],2'b0})+$signed(-{in[68],2'b0})+$signed(-in[12])+$signed({in[38],1'b0})+$signed(in[38])+$signed(sharing5_r)+$signed(1);
assign weighted_sum[175] = $signed({in[40],1'b0})+$signed(in[40])+$signed(-{in[42],2'b0})+$signed({in[68],1'b0})+$signed(-{in[69],2'b0})+$signed(-{in[70],2'b0})+$signed(-in[14])+$signed(sharing148_r)+$signed(1);
assign weighted_sum[176] = $signed(-{in[72],2'b0})+$signed(-in[16])+$signed({in[42],1'b0})+$signed(in[42])+$signed(-{in[44],2'b0})+$signed({in[70],1'b0})+$signed(-{in[71],2'b0})+$signed(sharing6_r)+$signed(1);
assign weighted_sum[177] = $signed({in[72],1'b0})+$signed(-{in[73],2'b0})+$signed(-{in[74],2'b0})+$signed(-in[18])+$signed({in[44],1'b0})+$signed(in[44])+$signed(-{in[46],2'b0})+$signed(sharing7_r)+$signed(1);
assign weighted_sum[178] = $signed(-{in[48],2'b0})+$signed({in[74],1'b0})+$signed(-{in[75],2'b0})+$signed(-{in[76],2'b0})+$signed(-in[20])+$signed({in[46],1'b0})+$signed(in[46])+$signed(sharing8_r)+$signed(1);
assign weighted_sum[179] = $signed({in[48],1'b0})+$signed(in[48])+$signed(-{in[50],2'b0})+$signed({in[76],1'b0})+$signed(-{in[77],2'b0})+$signed(-{in[78],2'b0})+$signed(-in[22])+$signed(sharing9_r)+$signed(1);
assign weighted_sum[180] = $signed(-{in[80],2'b0})+$signed(-in[24])+$signed({in[50],1'b0})+$signed(in[50])+$signed(-{in[52],2'b0})+$signed({in[78],1'b0})+$signed(-{in[79],2'b0})+$signed(sharing10_r)+$signed(1);
assign weighted_sum[181] = $signed({in[80],1'b0})+$signed(-{in[81],2'b0})+$signed(-{in[82],2'b0})+$signed(-in[26])+$signed({in[52],1'b0})+$signed(in[52])+$signed(-{in[54],2'b0})+$signed(sharing11_r)+$signed(1);
assign weighted_sum[182] = $signed({in[112],1'b0})+$signed(-{in[113],2'b0})+$signed(-{in[114],2'b0})+$signed(-in[58])+$signed({in[84],1'b0})+$signed(in[84])+$signed(-{in[86],2'b0})+$signed(sharing12_r)+$signed(1);
assign weighted_sum[183] = $signed(-{in[88],2'b0})+$signed({in[114],1'b0})+$signed(-{in[115],2'b0})+$signed(-{in[116],2'b0})+$signed(-in[60])+$signed({in[86],1'b0})+$signed(in[86])+$signed(sharing149_r)+$signed(1);
assign weighted_sum[184] = $signed({in[88],1'b0})+$signed(in[88])+$signed(-{in[90],2'b0})+$signed({in[116],1'b0})+$signed(-{in[117],2'b0})+$signed(-{in[118],2'b0})+$signed(-in[62])+$signed(sharing13_r)+$signed(1);
assign weighted_sum[185] = $signed(-{in[120],2'b0})+$signed(-in[64])+$signed({in[90],1'b0})+$signed(in[90])+$signed(-{in[92],2'b0})+$signed({in[118],1'b0})+$signed(-{in[119],2'b0})+$signed(sharing14_r)+$signed(1);
assign weighted_sum[186] = $signed({in[120],1'b0})+$signed(-{in[121],2'b0})+$signed(-{in[122],2'b0})+$signed(-in[66])+$signed({in[92],1'b0})+$signed(in[92])+$signed(-{in[94],2'b0})+$signed(sharing15_r)+$signed(1);
assign weighted_sum[187] = $signed(-{in[96],2'b0})+$signed({in[122],1'b0})+$signed(-{in[123],2'b0})+$signed(-{in[124],2'b0})+$signed(-in[68])+$signed({in[94],1'b0})+$signed(in[94])+$signed(sharing16_r)+$signed(1);
assign weighted_sum[188] = $signed({in[96],1'b0})+$signed(in[96])+$signed(-{in[98],2'b0})+$signed({in[124],1'b0})+$signed(-{in[125],2'b0})+$signed(-{in[126],2'b0})+$signed(-in[70])+$signed(sharing17_r)+$signed(1);
assign weighted_sum[189] = $signed(-{in[128],2'b0})+$signed(-in[72])+$signed({in[98],1'b0})+$signed(in[98])+$signed(-{in[100],2'b0})+$signed({in[126],1'b0})+$signed(-{in[127],2'b0})+$signed(sharing18_r)+$signed(1);
assign weighted_sum[190] = $signed({in[128],1'b0})+$signed(-{in[129],2'b0})+$signed(-{in[130],2'b0})+$signed(-in[74])+$signed({in[100],1'b0})+$signed(in[100])+$signed(-{in[102],2'b0})+$signed(sharing19_r)+$signed(1);
assign weighted_sum[191] = $signed(-{in[104],2'b0})+$signed({in[130],1'b0})+$signed(-{in[131],2'b0})+$signed(-{in[132],2'b0})+$signed(-in[76])+$signed({in[102],1'b0})+$signed(in[102])+$signed(sharing150_r)+$signed(1);
assign weighted_sum[192] = $signed({in[104],1'b0})+$signed(in[104])+$signed(-{in[106],2'b0})+$signed({in[132],1'b0})+$signed(-{in[133],2'b0})+$signed(-{in[134],2'b0})+$signed(-in[78])+$signed(sharing20_r)+$signed(1);
assign weighted_sum[193] = $signed(-{in[136],2'b0})+$signed(-in[80])+$signed({in[106],1'b0})+$signed(in[106])+$signed(-{in[108],2'b0})+$signed({in[134],1'b0})+$signed(-{in[135],2'b0})+$signed(sharing21_r)+$signed(1);
assign weighted_sum[194] = $signed({in[136],1'b0})+$signed(-{in[137],2'b0})+$signed(-{in[138],2'b0})+$signed(-in[82])+$signed({in[108],1'b0})+$signed(in[108])+$signed(-{in[110],2'b0})+$signed(sharing22_r)+$signed(1);
assign weighted_sum[195] = $signed({in[168],1'b0})+$signed(-{in[169],2'b0})+$signed(-{in[170],2'b0})+$signed(-in[114])+$signed({in[140],1'b0})+$signed(in[140])+$signed(-{in[142],2'b0})+$signed(sharing23_r)+$signed(1);
assign weighted_sum[196] = $signed(-{in[144],2'b0})+$signed({in[170],1'b0})+$signed(-{in[171],2'b0})+$signed(-{in[172],2'b0})+$signed(-in[116])+$signed({in[142],1'b0})+$signed(in[142])+$signed(sharing24_r)+$signed(1);
assign weighted_sum[197] = $signed({in[144],1'b0})+$signed(in[144])+$signed(-{in[146],2'b0})+$signed({in[172],1'b0})+$signed(-{in[173],2'b0})+$signed(-{in[174],2'b0})+$signed(-in[118])+$signed(sharing25_r)+$signed(1);
assign weighted_sum[198] = $signed(-{in[176],2'b0})+$signed(-in[120])+$signed({in[146],1'b0})+$signed(in[146])+$signed(-{in[148],2'b0})+$signed({in[174],1'b0})+$signed(-{in[175],2'b0})+$signed(sharing26_r)+$signed(1);
assign weighted_sum[199] = $signed({in[176],1'b0})+$signed(-{in[177],2'b0})+$signed(-{in[178],2'b0})+$signed(-in[122])+$signed({in[148],1'b0})+$signed(in[148])+$signed(-{in[150],2'b0})+$signed(sharing151_r)+$signed(1);
assign weighted_sum[200] = $signed(-{in[152],2'b0})+$signed({in[178],1'b0})+$signed(-{in[179],2'b0})+$signed(-{in[180],2'b0})+$signed(-in[124])+$signed({in[150],1'b0})+$signed(in[150])+$signed(sharing27_r)+$signed(1);
assign weighted_sum[201] = $signed({in[152],1'b0})+$signed(in[152])+$signed(-{in[154],2'b0})+$signed({in[180],1'b0})+$signed(-{in[181],2'b0})+$signed(-{in[182],2'b0})+$signed(-in[126])+$signed(sharing28_r)+$signed(1);
assign weighted_sum[202] = $signed(-{in[184],2'b0})+$signed(-in[128])+$signed({in[154],1'b0})+$signed(in[154])+$signed(-{in[156],2'b0})+$signed({in[182],1'b0})+$signed(-{in[183],2'b0})+$signed(sharing29_r)+$signed(1);
assign weighted_sum[203] = $signed({in[184],1'b0})+$signed(-{in[185],2'b0})+$signed(-{in[186],2'b0})+$signed(-in[130])+$signed({in[156],1'b0})+$signed(in[156])+$signed(-{in[158],2'b0})+$signed(sharing30_r)+$signed(1);
assign weighted_sum[204] = $signed(-{in[160],2'b0})+$signed({in[186],1'b0})+$signed(-{in[187],2'b0})+$signed(-{in[188],2'b0})+$signed(-in[132])+$signed({in[158],1'b0})+$signed(in[158])+$signed(sharing31_r)+$signed(1);
assign weighted_sum[205] = $signed({in[160],1'b0})+$signed(in[160])+$signed(-{in[162],2'b0})+$signed({in[188],1'b0})+$signed(-{in[189],2'b0})+$signed(-{in[190],2'b0})+$signed(-in[134])+$signed(sharing32_r)+$signed(1);
assign weighted_sum[206] = $signed(-{in[192],2'b0})+$signed(-in[136])+$signed({in[162],1'b0})+$signed(in[162])+$signed(-{in[164],2'b0})+$signed({in[190],1'b0})+$signed(-{in[191],2'b0})+$signed(sharing33_r)+$signed(1);
assign weighted_sum[207] = $signed({in[192],1'b0})+$signed(-{in[193],2'b0})+$signed(-{in[194],2'b0})+$signed(-in[138])+$signed({in[164],1'b0})+$signed(in[164])+$signed(-{in[166],2'b0})+$signed(sharing152_r)+$signed(1);
assign weighted_sum[208] = $signed({in[224],1'b0})+$signed(-{in[225],2'b0})+$signed(-{in[226],2'b0})+$signed(-in[170])+$signed({in[196],1'b0})+$signed(in[196])+$signed(-{in[198],2'b0})+$signed(sharing34_r)+$signed(1);
assign weighted_sum[209] = $signed(-{in[200],2'b0})+$signed({in[226],1'b0})+$signed(-{in[227],2'b0})+$signed(-{in[228],2'b0})+$signed(-in[172])+$signed({in[198],1'b0})+$signed(in[198])+$signed(sharing35_r)+$signed(1);
assign weighted_sum[210] = $signed({in[200],1'b0})+$signed(in[200])+$signed(-{in[202],2'b0})+$signed({in[228],1'b0})+$signed(-{in[229],2'b0})+$signed(-{in[230],2'b0})+$signed(-in[174])+$signed(sharing36_r)+$signed(1);
assign weighted_sum[211] = $signed(-{in[232],2'b0})+$signed(-in[176])+$signed({in[202],1'b0})+$signed(in[202])+$signed(-{in[204],2'b0})+$signed({in[230],1'b0})+$signed(-{in[231],2'b0})+$signed(sharing37_r)+$signed(1);
assign weighted_sum[212] = $signed({in[232],1'b0})+$signed(-{in[233],2'b0})+$signed(-{in[234],2'b0})+$signed(-in[178])+$signed({in[204],1'b0})+$signed(in[204])+$signed(-{in[206],2'b0})+$signed(sharing38_r)+$signed(1);
assign weighted_sum[213] = $signed(-{in[208],2'b0})+$signed({in[234],1'b0})+$signed(-{in[235],2'b0})+$signed(-{in[236],2'b0})+$signed(-in[180])+$signed({in[206],1'b0})+$signed(in[206])+$signed(sharing39_r)+$signed(1);
assign weighted_sum[214] = $signed({in[208],1'b0})+$signed(in[208])+$signed(-{in[210],2'b0})+$signed({in[236],1'b0})+$signed(-{in[237],2'b0})+$signed(-{in[238],2'b0})+$signed(-in[182])+$signed(sharing40_r)+$signed(1);
assign weighted_sum[215] = $signed(-{in[240],2'b0})+$signed(-in[184])+$signed({in[210],1'b0})+$signed(in[210])+$signed(-{in[212],2'b0})+$signed({in[238],1'b0})+$signed(-{in[239],2'b0})+$signed(sharing153_r)+$signed(1);
assign weighted_sum[216] = $signed({in[240],1'b0})+$signed(-{in[241],2'b0})+$signed(-{in[242],2'b0})+$signed(-in[186])+$signed({in[212],1'b0})+$signed(in[212])+$signed(-{in[214],2'b0})+$signed(sharing41_r)+$signed(1);
assign weighted_sum[217] = $signed(-{in[216],2'b0})+$signed({in[242],1'b0})+$signed(-{in[243],2'b0})+$signed(-{in[244],2'b0})+$signed(-in[188])+$signed({in[214],1'b0})+$signed(in[214])+$signed(sharing42_r)+$signed(1);
assign weighted_sum[218] = $signed({in[216],1'b0})+$signed(in[216])+$signed(-{in[218],2'b0})+$signed({in[244],1'b0})+$signed(-{in[245],2'b0})+$signed(-{in[246],2'b0})+$signed(-in[190])+$signed(sharing43_r)+$signed(1);
assign weighted_sum[219] = $signed(-{in[248],2'b0})+$signed(-in[192])+$signed({in[218],1'b0})+$signed(in[218])+$signed(-{in[220],2'b0})+$signed({in[246],1'b0})+$signed(-{in[247],2'b0})+$signed(sharing44_r)+$signed(1);
assign weighted_sum[220] = $signed({in[248],1'b0})+$signed(-{in[249],2'b0})+$signed(-{in[250],2'b0})+$signed(-in[194])+$signed({in[220],1'b0})+$signed(in[220])+$signed(-{in[222],2'b0})+$signed(sharing45_r)+$signed(1);
assign weighted_sum[221] = $signed({in[280],1'b0})+$signed(-{in[281],2'b0})+$signed(-{in[282],2'b0})+$signed(-in[226])+$signed({in[252],1'b0})+$signed(in[252])+$signed(-{in[254],2'b0})+$signed(sharing46_r)+$signed(1);
assign weighted_sum[222] = $signed(-{in[256],2'b0})+$signed({in[282],1'b0})+$signed(-{in[283],2'b0})+$signed(-{in[284],2'b0})+$signed(-in[228])+$signed({in[254],1'b0})+$signed(in[254])+$signed(sharing47_r)+$signed(1);
assign weighted_sum[223] = $signed({in[256],1'b0})+$signed(in[256])+$signed(-{in[258],2'b0})+$signed({in[284],1'b0})+$signed(-{in[285],2'b0})+$signed(-{in[286],2'b0})+$signed(-in[230])+$signed(sharing154_r)+$signed(1);
assign weighted_sum[224] = $signed(-{in[288],2'b0})+$signed(-in[232])+$signed({in[258],1'b0})+$signed(in[258])+$signed(-{in[260],2'b0})+$signed({in[286],1'b0})+$signed(-{in[287],2'b0})+$signed(sharing48_r)+$signed(1);
assign weighted_sum[225] = $signed({in[288],1'b0})+$signed(-{in[289],2'b0})+$signed(-{in[290],2'b0})+$signed(-in[234])+$signed({in[260],1'b0})+$signed(in[260])+$signed(-{in[262],2'b0})+$signed(sharing49_r)+$signed(1);
assign weighted_sum[226] = $signed(-{in[264],2'b0})+$signed({in[290],1'b0})+$signed(-{in[291],2'b0})+$signed(-{in[292],2'b0})+$signed(-in[236])+$signed({in[262],1'b0})+$signed(in[262])+$signed(sharing50_r)+$signed(1);
assign weighted_sum[227] = $signed({in[264],1'b0})+$signed(in[264])+$signed(-{in[266],2'b0})+$signed({in[292],1'b0})+$signed(-{in[293],2'b0})+$signed(-{in[294],2'b0})+$signed(-in[238])+$signed(sharing51_r)+$signed(1);
assign weighted_sum[228] = $signed(-{in[296],2'b0})+$signed(-in[240])+$signed({in[266],1'b0})+$signed(in[266])+$signed(-{in[268],2'b0})+$signed({in[294],1'b0})+$signed(-{in[295],2'b0})+$signed(sharing52_r)+$signed(1);
assign weighted_sum[229] = $signed({in[296],1'b0})+$signed(-{in[297],2'b0})+$signed(-{in[298],2'b0})+$signed(-in[242])+$signed({in[268],1'b0})+$signed(in[268])+$signed(-{in[270],2'b0})+$signed(sharing53_r)+$signed(1);
assign weighted_sum[230] = $signed(-{in[272],2'b0})+$signed({in[298],1'b0})+$signed(-{in[299],2'b0})+$signed(-{in[300],2'b0})+$signed(-in[244])+$signed({in[270],1'b0})+$signed(in[270])+$signed(sharing54_r)+$signed(1);
assign weighted_sum[231] = $signed({in[272],1'b0})+$signed(in[272])+$signed(-{in[274],2'b0})+$signed({in[300],1'b0})+$signed(-{in[301],2'b0})+$signed(-{in[302],2'b0})+$signed(-in[246])+$signed(sharing155_r)+$signed(1);
assign weighted_sum[232] = $signed(-{in[304],2'b0})+$signed(-in[248])+$signed({in[274],1'b0})+$signed(in[274])+$signed(-{in[276],2'b0})+$signed({in[302],1'b0})+$signed(-{in[303],2'b0})+$signed(sharing55_r)+$signed(1);
assign weighted_sum[233] = $signed({in[304],1'b0})+$signed(-{in[305],2'b0})+$signed(-{in[306],2'b0})+$signed(-in[250])+$signed({in[276],1'b0})+$signed(in[276])+$signed(-{in[278],2'b0})+$signed(sharing56_r)+$signed(1);
assign weighted_sum[234] = $signed({in[336],1'b0})+$signed(-{in[337],2'b0})+$signed(-{in[338],2'b0})+$signed(-in[282])+$signed({in[308],1'b0})+$signed(in[308])+$signed(-{in[310],2'b0})+$signed(sharing57_r)+$signed(1);
assign weighted_sum[235] = $signed(-{in[312],2'b0})+$signed({in[338],1'b0})+$signed(-{in[339],2'b0})+$signed(-{in[340],2'b0})+$signed(-in[284])+$signed({in[310],1'b0})+$signed(in[310])+$signed(sharing58_r)+$signed(1);
assign weighted_sum[236] = $signed({in[312],1'b0})+$signed(in[312])+$signed(-{in[314],2'b0})+$signed({in[340],1'b0})+$signed(-{in[341],2'b0})+$signed(-{in[342],2'b0})+$signed(-in[286])+$signed(sharing59_r)+$signed(1);
assign weighted_sum[237] = $signed(-{in[344],2'b0})+$signed(-in[288])+$signed({in[314],1'b0})+$signed(in[314])+$signed(-{in[316],2'b0})+$signed({in[342],1'b0})+$signed(-{in[343],2'b0})+$signed(sharing60_r)+$signed(1);
assign weighted_sum[238] = $signed({in[344],1'b0})+$signed(-{in[345],2'b0})+$signed(-{in[346],2'b0})+$signed(-in[290])+$signed({in[316],1'b0})+$signed(in[316])+$signed(-{in[318],2'b0})+$signed(sharing61_r)+$signed(1);
assign weighted_sum[239] = $signed(-{in[320],2'b0})+$signed({in[346],1'b0})+$signed(-{in[347],2'b0})+$signed(-{in[348],2'b0})+$signed(-in[292])+$signed({in[318],1'b0})+$signed(in[318])+$signed(sharing156_r)+$signed(1);
assign weighted_sum[240] = $signed({in[320],1'b0})+$signed(in[320])+$signed(-{in[322],2'b0})+$signed({in[348],1'b0})+$signed(-{in[349],2'b0})+$signed(-{in[350],2'b0})+$signed(-in[294])+$signed(sharing62_r)+$signed(1);
assign weighted_sum[241] = $signed(-{in[352],2'b0})+$signed(-in[296])+$signed({in[322],1'b0})+$signed(in[322])+$signed(-{in[324],2'b0})+$signed({in[350],1'b0})+$signed(-{in[351],2'b0})+$signed(sharing63_r)+$signed(1);
assign weighted_sum[242] = $signed({in[352],1'b0})+$signed(-{in[353],2'b0})+$signed(-{in[354],2'b0})+$signed(-in[298])+$signed({in[324],1'b0})+$signed(in[324])+$signed(-{in[326],2'b0})+$signed(sharing64_r)+$signed(1);
assign weighted_sum[243] = $signed(-{in[328],2'b0})+$signed({in[354],1'b0})+$signed(-{in[355],2'b0})+$signed(-{in[356],2'b0})+$signed(-in[300])+$signed({in[326],1'b0})+$signed(in[326])+$signed(sharing65_r)+$signed(1);
assign weighted_sum[244] = $signed({in[328],1'b0})+$signed(in[328])+$signed(-{in[330],2'b0})+$signed({in[356],1'b0})+$signed(-{in[357],2'b0})+$signed(-{in[358],2'b0})+$signed(-in[302])+$signed(sharing66_r)+$signed(1);
assign weighted_sum[245] = $signed(-{in[360],2'b0})+$signed(-in[304])+$signed({in[330],1'b0})+$signed(in[330])+$signed(-{in[332],2'b0})+$signed({in[358],1'b0})+$signed(-{in[359],2'b0})+$signed(sharing67_r)+$signed(1);
assign weighted_sum[246] = $signed({in[360],1'b0})+$signed(-{in[361],2'b0})+$signed(-{in[362],2'b0})+$signed(-in[306])+$signed({in[332],1'b0})+$signed(in[332])+$signed(-{in[334],2'b0})+$signed(sharing68_r)+$signed(1);
assign weighted_sum[247] = $signed({in[392],1'b0})+$signed(-{in[393],2'b0})+$signed(-{in[394],2'b0})+$signed(-in[338])+$signed({in[364],1'b0})+$signed(in[364])+$signed(-{in[366],2'b0})+$signed(sharing157_r)+$signed(1);
assign weighted_sum[248] = $signed(-{in[368],2'b0})+$signed({in[394],1'b0})+$signed(-{in[395],2'b0})+$signed(-{in[396],2'b0})+$signed(-in[340])+$signed({in[366],1'b0})+$signed(in[366])+$signed(sharing69_r)+$signed(1);
assign weighted_sum[249] = $signed({in[368],1'b0})+$signed(in[368])+$signed(-{in[370],2'b0})+$signed({in[396],1'b0})+$signed(-{in[397],2'b0})+$signed(-{in[398],2'b0})+$signed(-in[342])+$signed(sharing70_r)+$signed(1);
assign weighted_sum[250] = $signed(-{in[400],2'b0})+$signed(-in[344])+$signed({in[370],1'b0})+$signed(in[370])+$signed(-{in[372],2'b0})+$signed({in[398],1'b0})+$signed(-{in[399],2'b0})+$signed(sharing71_r)+$signed(1);
assign weighted_sum[251] = $signed({in[400],1'b0})+$signed(-{in[401],2'b0})+$signed(-{in[402],2'b0})+$signed(-in[346])+$signed({in[372],1'b0})+$signed(in[372])+$signed(-{in[374],2'b0})+$signed(sharing72_r)+$signed(1);
assign weighted_sum[252] = $signed(-{in[376],2'b0})+$signed({in[402],1'b0})+$signed(-{in[403],2'b0})+$signed(-{in[404],2'b0})+$signed(-in[348])+$signed({in[374],1'b0})+$signed(in[374])+$signed(sharing73_r)+$signed(1);
assign weighted_sum[253] = $signed({in[376],1'b0})+$signed(in[376])+$signed(-{in[378],2'b0})+$signed({in[404],1'b0})+$signed(-{in[405],2'b0})+$signed(-{in[406],2'b0})+$signed(-in[350])+$signed(sharing74_r)+$signed(1);
assign weighted_sum[254] = $signed(-{in[408],2'b0})+$signed(-in[352])+$signed({in[378],1'b0})+$signed(in[378])+$signed(-{in[380],2'b0})+$signed({in[406],1'b0})+$signed(-{in[407],2'b0})+$signed(sharing75_r)+$signed(1);
assign weighted_sum[255] = $signed({in[408],1'b0})+$signed(-{in[409],2'b0})+$signed(-{in[410],2'b0})+$signed(-in[354])+$signed({in[380],1'b0})+$signed(in[380])+$signed(-{in[382],2'b0})+$signed(sharing158_r)+$signed(1);
assign weighted_sum[256] = $signed(-{in[384],2'b0})+$signed({in[410],1'b0})+$signed(-{in[411],2'b0})+$signed(-{in[412],2'b0})+$signed(-in[356])+$signed({in[382],1'b0})+$signed(in[382])+$signed(sharing76_r)+$signed(1);
assign weighted_sum[257] = $signed({in[384],1'b0})+$signed(in[384])+$signed(-{in[386],2'b0})+$signed({in[412],1'b0})+$signed(-{in[413],2'b0})+$signed(-{in[414],2'b0})+$signed(-in[358])+$signed(sharing77_r)+$signed(1);
assign weighted_sum[258] = $signed(-{in[416],2'b0})+$signed(-in[360])+$signed({in[386],1'b0})+$signed(in[386])+$signed(-{in[388],2'b0})+$signed({in[414],1'b0})+$signed(-{in[415],2'b0})+$signed(sharing78_r)+$signed(1);
assign weighted_sum[259] = $signed({in[416],1'b0})+$signed(-{in[417],2'b0})+$signed(-{in[418],2'b0})+$signed(-in[362])+$signed({in[388],1'b0})+$signed(in[388])+$signed(-{in[390],2'b0})+$signed(sharing79_r)+$signed(1);
assign weighted_sum[260] = $signed({in[448],1'b0})+$signed(-{in[449],2'b0})+$signed(-{in[450],2'b0})+$signed(-in[394])+$signed({in[420],1'b0})+$signed(in[420])+$signed(-{in[422],2'b0})+$signed(sharing80_r)+$signed(1);
assign weighted_sum[261] = $signed(-{in[424],2'b0})+$signed({in[450],1'b0})+$signed(-{in[451],2'b0})+$signed(-{in[452],2'b0})+$signed(-in[396])+$signed({in[422],1'b0})+$signed(in[422])+$signed(sharing81_r)+$signed(1);
assign weighted_sum[262] = $signed({in[424],1'b0})+$signed(in[424])+$signed(-{in[426],2'b0})+$signed({in[452],1'b0})+$signed(-{in[453],2'b0})+$signed(-{in[454],2'b0})+$signed(-in[398])+$signed(sharing82_r)+$signed(1);
assign weighted_sum[263] = $signed(-{in[456],2'b0})+$signed(-in[400])+$signed({in[426],1'b0})+$signed(in[426])+$signed(-{in[428],2'b0})+$signed({in[454],1'b0})+$signed(-{in[455],2'b0})+$signed(sharing159_r)+$signed(1);
assign weighted_sum[264] = $signed({in[456],1'b0})+$signed(-{in[457],2'b0})+$signed(-{in[458],2'b0})+$signed(-in[402])+$signed({in[428],1'b0})+$signed(in[428])+$signed(-{in[430],2'b0})+$signed(sharing83_r)+$signed(1);
assign weighted_sum[265] = $signed(-{in[432],2'b0})+$signed({in[458],1'b0})+$signed(-{in[459],2'b0})+$signed(-{in[460],2'b0})+$signed(-in[404])+$signed({in[430],1'b0})+$signed(in[430])+$signed(sharing84_r)+$signed(1);
assign weighted_sum[266] = $signed({in[432],1'b0})+$signed(in[432])+$signed(-{in[434],2'b0})+$signed({in[460],1'b0})+$signed(-{in[461],2'b0})+$signed(-{in[462],2'b0})+$signed(-in[406])+$signed(sharing85_r)+$signed(1);
assign weighted_sum[267] = $signed(-{in[464],2'b0})+$signed(-in[408])+$signed({in[434],1'b0})+$signed(in[434])+$signed(-{in[436],2'b0})+$signed({in[462],1'b0})+$signed(-{in[463],2'b0})+$signed(sharing86_r)+$signed(1);
assign weighted_sum[268] = $signed({in[464],1'b0})+$signed(-{in[465],2'b0})+$signed(-{in[466],2'b0})+$signed(-in[410])+$signed({in[436],1'b0})+$signed(in[436])+$signed(-{in[438],2'b0})+$signed(sharing87_r)+$signed(1);
assign weighted_sum[269] = $signed(-{in[440],2'b0})+$signed({in[466],1'b0})+$signed(-{in[467],2'b0})+$signed(-{in[468],2'b0})+$signed(-in[412])+$signed({in[438],1'b0})+$signed(in[438])+$signed(sharing88_r)+$signed(1);
assign weighted_sum[270] = $signed({in[440],1'b0})+$signed(in[440])+$signed(-{in[442],2'b0})+$signed({in[468],1'b0})+$signed(-{in[469],2'b0})+$signed(-{in[470],2'b0})+$signed(-in[414])+$signed(sharing89_r)+$signed(1);
assign weighted_sum[271] = $signed(-{in[472],2'b0})+$signed(-in[416])+$signed({in[442],1'b0})+$signed(in[442])+$signed(-{in[444],2'b0})+$signed({in[470],1'b0})+$signed(-{in[471],2'b0})+$signed(sharing160_r)+$signed(1);
assign weighted_sum[272] = $signed({in[472],1'b0})+$signed(-{in[473],2'b0})+$signed(-{in[474],2'b0})+$signed(-in[418])+$signed({in[444],1'b0})+$signed(in[444])+$signed(-{in[446],2'b0})+$signed(sharing90_r)+$signed(1);
assign weighted_sum[273] = $signed({in[504],1'b0})+$signed(-{in[505],2'b0})+$signed(-{in[506],2'b0})+$signed(-in[450])+$signed({in[476],1'b0})+$signed(in[476])+$signed(-{in[478],2'b0})+$signed(sharing91_r)+$signed(1);
assign weighted_sum[274] = $signed(-{in[480],2'b0})+$signed({in[506],1'b0})+$signed(-{in[507],2'b0})+$signed(-{in[508],2'b0})+$signed(-in[452])+$signed({in[478],1'b0})+$signed(in[478])+$signed(sharing92_r)+$signed(1);
assign weighted_sum[275] = $signed({in[480],1'b0})+$signed(in[480])+$signed(-{in[482],2'b0})+$signed({in[508],1'b0})+$signed(-{in[509],2'b0})+$signed(-{in[510],2'b0})+$signed(-in[454])+$signed(sharing93_r)+$signed(1);
assign weighted_sum[276] = $signed(-{in[512],2'b0})+$signed(-in[456])+$signed({in[482],1'b0})+$signed(in[482])+$signed(-{in[484],2'b0})+$signed({in[510],1'b0})+$signed(-{in[511],2'b0})+$signed(sharing94_r)+$signed(1);
assign weighted_sum[277] = $signed({in[512],1'b0})+$signed(-{in[513],2'b0})+$signed(-{in[514],2'b0})+$signed(-in[458])+$signed({in[484],1'b0})+$signed(in[484])+$signed(-{in[486],2'b0})+$signed(sharing95_r)+$signed(1);
assign weighted_sum[278] = $signed(-{in[488],2'b0})+$signed({in[514],1'b0})+$signed(-{in[515],2'b0})+$signed(-{in[516],2'b0})+$signed(-in[460])+$signed({in[486],1'b0})+$signed(in[486])+$signed(sharing96_r)+$signed(1);
assign weighted_sum[279] = $signed({in[488],1'b0})+$signed(in[488])+$signed(-{in[490],2'b0})+$signed({in[516],1'b0})+$signed(-{in[517],2'b0})+$signed(-{in[518],2'b0})+$signed(-in[462])+$signed(sharing161_r)+$signed(1);
assign weighted_sum[280] = $signed(-{in[520],2'b0})+$signed(-in[464])+$signed({in[490],1'b0})+$signed(in[490])+$signed(-{in[492],2'b0})+$signed({in[518],1'b0})+$signed(-{in[519],2'b0})+$signed(sharing97_r)+$signed(1);
assign weighted_sum[281] = $signed({in[520],1'b0})+$signed(-{in[521],2'b0})+$signed(-{in[522],2'b0})+$signed(-in[466])+$signed({in[492],1'b0})+$signed(in[492])+$signed(-{in[494],2'b0})+$signed(sharing98_r)+$signed(1);
assign weighted_sum[282] = $signed(-{in[496],2'b0})+$signed({in[522],1'b0})+$signed(-{in[523],2'b0})+$signed(-{in[524],2'b0})+$signed(-in[468])+$signed({in[494],1'b0})+$signed(in[494])+$signed(sharing99_r)+$signed(1);
assign weighted_sum[283] = $signed({in[496],1'b0})+$signed(in[496])+$signed(-{in[498],2'b0})+$signed({in[524],1'b0})+$signed(-{in[525],2'b0})+$signed(-{in[526],2'b0})+$signed(-in[470])+$signed(sharing100_r)+$signed(1);
assign weighted_sum[284] = $signed(-{in[528],2'b0})+$signed(-in[472])+$signed({in[498],1'b0})+$signed(in[498])+$signed(-{in[500],2'b0})+$signed({in[526],1'b0})+$signed(-{in[527],2'b0})+$signed(sharing101_r)+$signed(1);
assign weighted_sum[285] = $signed({in[528],1'b0})+$signed(-{in[529],2'b0})+$signed(-{in[530],2'b0})+$signed(-in[474])+$signed({in[500],1'b0})+$signed(in[500])+$signed(-{in[502],2'b0})+$signed(sharing102_r)+$signed(1);
assign weighted_sum[286] = $signed({in[560],1'b0})+$signed(-{in[561],2'b0})+$signed(-{in[562],2'b0})+$signed(-in[506])+$signed({in[532],1'b0})+$signed(in[532])+$signed(-{in[534],2'b0})+$signed(sharing103_r)+$signed(1);
assign weighted_sum[287] = $signed(-{in[536],2'b0})+$signed({in[562],1'b0})+$signed(-{in[563],2'b0})+$signed(-{in[564],2'b0})+$signed(-in[508])+$signed({in[534],1'b0})+$signed(in[534])+$signed(sharing162_r)+$signed(1);
assign weighted_sum[288] = $signed({in[536],1'b0})+$signed(in[536])+$signed(-{in[538],2'b0})+$signed({in[564],1'b0})+$signed(-{in[565],2'b0})+$signed(-{in[566],2'b0})+$signed(-in[510])+$signed(sharing104_r)+$signed(1);
assign weighted_sum[289] = $signed(-{in[568],2'b0})+$signed(-in[512])+$signed({in[538],1'b0})+$signed(in[538])+$signed(-{in[540],2'b0})+$signed({in[566],1'b0})+$signed(-{in[567],2'b0})+$signed(sharing105_r)+$signed(1);
assign weighted_sum[290] = $signed({in[568],1'b0})+$signed(-{in[569],2'b0})+$signed(-{in[570],2'b0})+$signed(-in[514])+$signed({in[540],1'b0})+$signed(in[540])+$signed(-{in[542],2'b0})+$signed(sharing106_r)+$signed(1);
assign weighted_sum[291] = $signed(-{in[544],2'b0})+$signed({in[570],1'b0})+$signed(-{in[571],2'b0})+$signed(-{in[572],2'b0})+$signed(-in[516])+$signed({in[542],1'b0})+$signed(in[542])+$signed(sharing107_r)+$signed(1);
assign weighted_sum[292] = $signed({in[544],1'b0})+$signed(in[544])+$signed(-{in[546],2'b0})+$signed({in[572],1'b0})+$signed(-{in[573],2'b0})+$signed(-{in[574],2'b0})+$signed(-in[518])+$signed(sharing108_r)+$signed(1);
assign weighted_sum[293] = $signed(-{in[576],2'b0})+$signed(-in[520])+$signed({in[546],1'b0})+$signed(in[546])+$signed(-{in[548],2'b0})+$signed({in[574],1'b0})+$signed(-{in[575],2'b0})+$signed(sharing109_r)+$signed(1);
assign weighted_sum[294] = $signed({in[576],1'b0})+$signed(-{in[577],2'b0})+$signed(-{in[578],2'b0})+$signed(-in[522])+$signed({in[548],1'b0})+$signed(in[548])+$signed(-{in[550],2'b0})+$signed(sharing110_r)+$signed(1);
assign weighted_sum[295] = $signed(-{in[552],2'b0})+$signed({in[578],1'b0})+$signed(-{in[579],2'b0})+$signed(-{in[580],2'b0})+$signed(-in[524])+$signed({in[550],1'b0})+$signed(in[550])+$signed(sharing163_r)+$signed(1);
assign weighted_sum[296] = $signed({in[552],1'b0})+$signed(in[552])+$signed(-{in[554],2'b0})+$signed({in[580],1'b0})+$signed(-{in[581],2'b0})+$signed(-{in[582],2'b0})+$signed(-in[526])+$signed(sharing111_r)+$signed(1);
assign weighted_sum[297] = $signed(-{in[584],2'b0})+$signed(-in[528])+$signed({in[554],1'b0})+$signed(in[554])+$signed(-{in[556],2'b0})+$signed({in[582],1'b0})+$signed(-{in[583],2'b0})+$signed(sharing112_r)+$signed(1);
assign weighted_sum[298] = $signed({in[584],1'b0})+$signed(-{in[585],2'b0})+$signed(-{in[586],2'b0})+$signed(-in[530])+$signed({in[556],1'b0})+$signed(in[556])+$signed(-{in[558],2'b0})+$signed(sharing113_r)+$signed(1);
assign weighted_sum[299] = $signed({in[616],1'b0})+$signed(-{in[617],2'b0})+$signed(-{in[618],2'b0})+$signed(-in[562])+$signed({in[588],1'b0})+$signed(in[588])+$signed(-{in[590],2'b0})+$signed(sharing114_r)+$signed(1);
assign weighted_sum[300] = $signed(-{in[592],2'b0})+$signed({in[618],1'b0})+$signed(-{in[619],2'b0})+$signed(-{in[620],2'b0})+$signed(-in[564])+$signed({in[590],1'b0})+$signed(in[590])+$signed(sharing115_r)+$signed(1);
assign weighted_sum[301] = $signed({in[592],1'b0})+$signed(in[592])+$signed(-{in[594],2'b0})+$signed({in[620],1'b0})+$signed(-{in[621],2'b0})+$signed(-{in[622],2'b0})+$signed(-in[566])+$signed(sharing116_r)+$signed(1);
assign weighted_sum[302] = $signed(-{in[624],2'b0})+$signed(-in[568])+$signed({in[594],1'b0})+$signed(in[594])+$signed(-{in[596],2'b0})+$signed({in[622],1'b0})+$signed(-{in[623],2'b0})+$signed(sharing117_r)+$signed(1);
assign weighted_sum[303] = $signed({in[624],1'b0})+$signed(-{in[625],2'b0})+$signed(-{in[626],2'b0})+$signed(-in[570])+$signed({in[596],1'b0})+$signed(in[596])+$signed(-{in[598],2'b0})+$signed(sharing164_r)+$signed(1);
assign weighted_sum[304] = $signed(-{in[600],2'b0})+$signed({in[626],1'b0})+$signed(-{in[627],2'b0})+$signed(-{in[628],2'b0})+$signed(-in[572])+$signed({in[598],1'b0})+$signed(in[598])+$signed(sharing118_r)+$signed(1);
assign weighted_sum[305] = $signed({in[600],1'b0})+$signed(in[600])+$signed(-{in[602],2'b0})+$signed({in[628],1'b0})+$signed(-{in[629],2'b0})+$signed(-{in[630],2'b0})+$signed(-in[574])+$signed(sharing119_r)+$signed(1);
assign weighted_sum[306] = $signed(-{in[632],2'b0})+$signed(-in[576])+$signed({in[602],1'b0})+$signed(in[602])+$signed(-{in[604],2'b0})+$signed({in[630],1'b0})+$signed(-{in[631],2'b0})+$signed(sharing120_r)+$signed(1);
assign weighted_sum[307] = $signed({in[632],1'b0})+$signed(-{in[633],2'b0})+$signed(-{in[634],2'b0})+$signed(-in[578])+$signed({in[604],1'b0})+$signed(in[604])+$signed(-{in[606],2'b0})+$signed(sharing121_r)+$signed(1);
assign weighted_sum[308] = $signed(-{in[608],2'b0})+$signed({in[634],1'b0})+$signed(-{in[635],2'b0})+$signed(-{in[636],2'b0})+$signed(-in[580])+$signed({in[606],1'b0})+$signed(in[606])+$signed(sharing122_r)+$signed(1);
assign weighted_sum[309] = $signed({in[608],1'b0})+$signed(in[608])+$signed(-{in[610],2'b0})+$signed({in[636],1'b0})+$signed(-{in[637],2'b0})+$signed(-{in[638],2'b0})+$signed(-in[582])+$signed(sharing123_r)+$signed(1);
assign weighted_sum[310] = $signed(-{in[640],2'b0})+$signed(-in[584])+$signed({in[610],1'b0})+$signed(in[610])+$signed(-{in[612],2'b0})+$signed({in[638],1'b0})+$signed(-{in[639],2'b0})+$signed(sharing124_r)+$signed(1);
assign weighted_sum[311] = $signed({in[640],1'b0})+$signed(-{in[641],2'b0})+$signed(-{in[642],2'b0})+$signed(-in[586])+$signed({in[612],1'b0})+$signed(in[612])+$signed(-{in[614],2'b0})+$signed(sharing165_r)+$signed(1);
assign weighted_sum[312] = $signed({in[672],1'b0})+$signed(-{in[673],2'b0})+$signed(-{in[674],2'b0})+$signed(-in[618])+$signed({in[644],1'b0})+$signed(in[644])+$signed(-{in[646],2'b0})+$signed(sharing125_r)+$signed(1);
assign weighted_sum[313] = $signed(-{in[648],2'b0})+$signed({in[674],1'b0})+$signed(-{in[675],2'b0})+$signed(-{in[676],2'b0})+$signed(-in[620])+$signed({in[646],1'b0})+$signed(in[646])+$signed(sharing126_r)+$signed(1);
assign weighted_sum[314] = $signed({in[648],1'b0})+$signed(in[648])+$signed(-{in[650],2'b0})+$signed({in[676],1'b0})+$signed(-{in[677],2'b0})+$signed(-{in[678],2'b0})+$signed(-in[622])+$signed(sharing127_r)+$signed(1);
assign weighted_sum[315] = $signed(-{in[680],2'b0})+$signed(-in[624])+$signed({in[650],1'b0})+$signed(in[650])+$signed(-{in[652],2'b0})+$signed({in[678],1'b0})+$signed(-{in[679],2'b0})+$signed(sharing128_r)+$signed(1);
assign weighted_sum[316] = $signed({in[680],1'b0})+$signed(-{in[681],2'b0})+$signed(-{in[682],2'b0})+$signed(-in[626])+$signed({in[652],1'b0})+$signed(in[652])+$signed(-{in[654],2'b0})+$signed(sharing129_r)+$signed(1);
assign weighted_sum[317] = $signed(-{in[656],2'b0})+$signed({in[682],1'b0})+$signed(-{in[683],2'b0})+$signed(-{in[684],2'b0})+$signed(-in[628])+$signed({in[654],1'b0})+$signed(in[654])+$signed(sharing130_r)+$signed(1);
assign weighted_sum[318] = $signed({in[656],1'b0})+$signed(in[656])+$signed(-{in[658],2'b0})+$signed({in[684],1'b0})+$signed(-{in[685],2'b0})+$signed(-{in[686],2'b0})+$signed(-in[630])+$signed(sharing131_r)+$signed(1);
assign weighted_sum[319] = $signed(-{in[688],2'b0})+$signed(-in[632])+$signed({in[658],1'b0})+$signed(in[658])+$signed(-{in[660],2'b0})+$signed({in[686],1'b0})+$signed(-{in[687],2'b0})+$signed(sharing166_r)+$signed(1);
assign weighted_sum[320] = $signed({in[688],1'b0})+$signed(-{in[689],2'b0})+$signed(-{in[690],2'b0})+$signed(-in[634])+$signed({in[660],1'b0})+$signed(in[660])+$signed(-{in[662],2'b0})+$signed(sharing132_r)+$signed(1);
assign weighted_sum[321] = $signed(-{in[664],2'b0})+$signed({in[690],1'b0})+$signed(-{in[691],2'b0})+$signed(-{in[692],2'b0})+$signed(-in[636])+$signed({in[662],1'b0})+$signed(in[662])+$signed(sharing133_r)+$signed(1);
assign weighted_sum[322] = $signed({in[664],1'b0})+$signed(in[664])+$signed(-{in[666],2'b0})+$signed({in[692],1'b0})+$signed(-{in[693],2'b0})+$signed(-{in[694],2'b0})+$signed(-in[638])+$signed(sharing134_r)+$signed(1);
assign weighted_sum[323] = $signed(-{in[696],2'b0})+$signed(-in[640])+$signed({in[666],1'b0})+$signed(in[666])+$signed(-{in[668],2'b0})+$signed({in[694],1'b0})+$signed(-{in[695],2'b0})+$signed(sharing135_r)+$signed(1);
assign weighted_sum[324] = $signed({in[696],1'b0})+$signed(-{in[697],2'b0})+$signed(-{in[698],2'b0})+$signed(-in[642])+$signed({in[668],1'b0})+$signed(in[668])+$signed(-{in[670],2'b0})+$signed(sharing136_r)+$signed(1);
assign weighted_sum[325] = $signed({in[728],1'b0})+$signed(-{in[729],2'b0})+$signed(-{in[730],2'b0})+$signed(-in[674])+$signed({in[700],1'b0})+$signed(in[700])+$signed(-{in[702],2'b0})+$signed(sharing137_r)+$signed(1);
assign weighted_sum[326] = $signed(-{in[704],2'b0})+$signed({in[730],1'b0})+$signed(-{in[731],2'b0})+$signed(-{in[732],2'b0})+$signed(-in[676])+$signed({in[702],1'b0})+$signed(in[702])+$signed(sharing138_r)+$signed(1);
assign weighted_sum[327] = $signed({in[704],1'b0})+$signed(in[704])+$signed(-{in[706],2'b0})+$signed({in[732],1'b0})+$signed(-{in[733],2'b0})+$signed(-{in[734],2'b0})+$signed(-in[678])+$signed(sharing167_r)+$signed(1);
assign weighted_sum[328] = $signed(-{in[736],2'b0})+$signed(-in[680])+$signed({in[706],1'b0})+$signed(in[706])+$signed(-{in[708],2'b0})+$signed({in[734],1'b0})+$signed(-{in[735],2'b0})+$signed(sharing139_r)+$signed(1);
assign weighted_sum[329] = $signed({in[736],1'b0})+$signed(-{in[737],2'b0})+$signed(-{in[738],2'b0})+$signed(-in[682])+$signed({in[708],1'b0})+$signed(in[708])+$signed(-{in[710],2'b0})+$signed(sharing140_r)+$signed(1);
assign weighted_sum[330] = $signed(-{in[712],2'b0})+$signed({in[738],1'b0})+$signed(-{in[739],2'b0})+$signed(-{in[740],2'b0})+$signed(-in[684])+$signed({in[710],1'b0})+$signed(in[710])+$signed(sharing141_r)+$signed(1);
assign weighted_sum[331] = $signed({in[712],1'b0})+$signed(in[712])+$signed(-{in[714],2'b0})+$signed({in[740],1'b0})+$signed(-{in[741],2'b0})+$signed(-{in[742],2'b0})+$signed(-in[686])+$signed(sharing142_r)+$signed(1);
assign weighted_sum[332] = $signed(-{in[744],2'b0})+$signed(-in[688])+$signed({in[714],1'b0})+$signed(in[714])+$signed(-{in[716],2'b0})+$signed({in[742],1'b0})+$signed(-{in[743],2'b0})+$signed(sharing143_r)+$signed(1);
assign weighted_sum[333] = $signed({in[744],1'b0})+$signed(-{in[745],2'b0})+$signed(-{in[746],2'b0})+$signed(-in[690])+$signed({in[716],1'b0})+$signed(in[716])+$signed(-{in[718],2'b0})+$signed(sharing144_r)+$signed(1);
assign weighted_sum[334] = $signed(-{in[720],2'b0})+$signed({in[746],1'b0})+$signed(-{in[747],2'b0})+$signed(-{in[748],2'b0})+$signed(-in[692])+$signed({in[718],1'b0})+$signed(in[718])+$signed(sharing145_r)+$signed(1);
assign weighted_sum[335] = $signed({in[720],1'b0})+$signed(in[720])+$signed(-{in[722],2'b0})+$signed({in[748],1'b0})+$signed(-{in[749],2'b0})+$signed(-{in[750],2'b0})+$signed(-in[694])+$signed(sharing168_r)+$signed(1);
assign weighted_sum[336] = $signed(-{in[752],2'b0})+$signed(-in[696])+$signed({in[722],1'b0})+$signed(in[722])+$signed(-{in[724],2'b0})+$signed({in[750],1'b0})+$signed(-{in[751],2'b0})+$signed(sharing146_r)+$signed(1);
assign weighted_sum[337] = $signed({in[752],1'b0})+$signed(-{in[753],2'b0})+$signed(-{in[754],2'b0})+$signed(-in[698])+$signed({in[724],1'b0})+$signed(in[724])+$signed(-{in[726],2'b0})+$signed(sharing147_r)+$signed(1);
assign weighted_sum[338] = $signed(-{in[56],3'b0})+$signed(-{in[57],3'b0})+$signed({in[1],1'b0})+$signed({in[2],2'b0})+$signed(-{in[58],1'b0})+$signed(in[2])+$signed(-{in[28],2'b0})+$signed({in[29],1'b0})+$signed({in[30],1'b0})+$signed(in[30])+$signed(sharing0_r)+$signed(-1);
assign weighted_sum[339] = $signed({in[32],1'b0})+$signed(in[32])+$signed(-{in[58],3'b0})+$signed(-{in[59],3'b0})+$signed({in[3],1'b0})+$signed({in[4],2'b0})+$signed(-{in[60],1'b0})+$signed(in[4])+$signed(-{in[30],2'b0})+$signed({in[31],1'b0})+$signed(sharing1_r)+$signed(-1);
assign weighted_sum[340] = $signed(-{in[32],2'b0})+$signed({in[33],1'b0})+$signed({in[34],1'b0})+$signed(in[34])+$signed(-{in[60],3'b0})+$signed(-{in[61],3'b0})+$signed({in[5],1'b0})+$signed({in[6],2'b0})+$signed(-{in[62],1'b0})+$signed(in[6])+$signed(sharing2_r)+$signed(-1);
assign weighted_sum[341] = $signed({in[8],2'b0})+$signed(-{in[64],1'b0})+$signed(in[8])+$signed(-{in[34],2'b0})+$signed({in[35],1'b0})+$signed({in[36],1'b0})+$signed(in[36])+$signed(-{in[62],3'b0})+$signed(-{in[63],3'b0})+$signed({in[7],1'b0})+$signed(sharing3_r)+$signed(-1);
assign weighted_sum[342] = $signed(-{in[64],3'b0})+$signed(-{in[65],3'b0})+$signed({in[9],1'b0})+$signed({in[10],2'b0})+$signed(-{in[66],1'b0})+$signed(in[10])+$signed(-{in[36],2'b0})+$signed({in[37],1'b0})+$signed({in[38],1'b0})+$signed(in[38])+$signed(sharing4_r)+$signed(-1);
assign weighted_sum[343] = $signed({in[40],1'b0})+$signed(in[40])+$signed(-{in[66],3'b0})+$signed(-{in[67],3'b0})+$signed({in[11],1'b0})+$signed({in[12],2'b0})+$signed(-{in[68],1'b0})+$signed(in[12])+$signed(-{in[38],2'b0})+$signed({in[39],1'b0})+$signed(sharing5_r)+$signed(-1);
assign weighted_sum[344] = $signed(-{in[40],2'b0})+$signed({in[41],1'b0})+$signed({in[42],1'b0})+$signed(in[42])+$signed(-{in[68],3'b0})+$signed(-{in[69],3'b0})+$signed({in[13],1'b0})+$signed({in[14],2'b0})+$signed(-{in[70],1'b0})+$signed(in[14])+$signed(sharing148_r)+$signed(-1);
assign weighted_sum[345] = $signed({in[16],2'b0})+$signed(-{in[72],1'b0})+$signed(in[16])+$signed(-{in[42],2'b0})+$signed({in[43],1'b0})+$signed({in[44],1'b0})+$signed(in[44])+$signed(-{in[70],3'b0})+$signed(-{in[71],3'b0})+$signed({in[15],1'b0})+$signed(sharing6_r)+$signed(-1);
assign weighted_sum[346] = $signed(-{in[72],3'b0})+$signed(-{in[73],3'b0})+$signed({in[17],1'b0})+$signed({in[18],2'b0})+$signed(-{in[74],1'b0})+$signed(in[18])+$signed(-{in[44],2'b0})+$signed({in[45],1'b0})+$signed({in[46],1'b0})+$signed(in[46])+$signed(sharing7_r)+$signed(-1);
assign weighted_sum[347] = $signed({in[48],1'b0})+$signed(in[48])+$signed(-{in[74],3'b0})+$signed(-{in[75],3'b0})+$signed({in[19],1'b0})+$signed({in[20],2'b0})+$signed(-{in[76],1'b0})+$signed(in[20])+$signed(-{in[46],2'b0})+$signed({in[47],1'b0})+$signed(sharing8_r)+$signed(-1);
assign weighted_sum[348] = $signed(-{in[48],2'b0})+$signed({in[49],1'b0})+$signed({in[50],1'b0})+$signed(in[50])+$signed(-{in[76],3'b0})+$signed(-{in[77],3'b0})+$signed({in[21],1'b0})+$signed({in[22],2'b0})+$signed(-{in[78],1'b0})+$signed(in[22])+$signed(sharing9_r)+$signed(-1);
assign weighted_sum[349] = $signed({in[24],2'b0})+$signed(-{in[80],1'b0})+$signed(in[24])+$signed(-{in[50],2'b0})+$signed({in[51],1'b0})+$signed({in[52],1'b0})+$signed(in[52])+$signed(-{in[78],3'b0})+$signed(-{in[79],3'b0})+$signed({in[23],1'b0})+$signed(sharing10_r)+$signed(-1);
assign weighted_sum[350] = $signed(-{in[80],3'b0})+$signed(-{in[81],3'b0})+$signed({in[25],1'b0})+$signed({in[26],2'b0})+$signed(-{in[82],1'b0})+$signed(in[26])+$signed(-{in[52],2'b0})+$signed({in[53],1'b0})+$signed({in[54],1'b0})+$signed(in[54])+$signed(sharing11_r)+$signed(-1);
assign weighted_sum[351] = $signed(-{in[112],3'b0})+$signed(-{in[113],3'b0})+$signed({in[57],1'b0})+$signed({in[58],2'b0})+$signed(-{in[114],1'b0})+$signed(in[58])+$signed(-{in[84],2'b0})+$signed({in[85],1'b0})+$signed({in[86],1'b0})+$signed(in[86])+$signed(sharing12_r)+$signed(-1);
assign weighted_sum[352] = $signed({in[88],1'b0})+$signed(in[88])+$signed(-{in[114],3'b0})+$signed(-{in[115],3'b0})+$signed({in[59],1'b0})+$signed({in[60],2'b0})+$signed(-{in[116],1'b0})+$signed(in[60])+$signed(-{in[86],2'b0})+$signed({in[87],1'b0})+$signed(sharing149_r)+$signed(-1);
assign weighted_sum[353] = $signed(-{in[88],2'b0})+$signed({in[89],1'b0})+$signed({in[90],1'b0})+$signed(in[90])+$signed(-{in[116],3'b0})+$signed(-{in[117],3'b0})+$signed({in[61],1'b0})+$signed({in[62],2'b0})+$signed(-{in[118],1'b0})+$signed(in[62])+$signed(sharing13_r)+$signed(-1);
assign weighted_sum[354] = $signed({in[64],2'b0})+$signed(-{in[120],1'b0})+$signed(in[64])+$signed(-{in[90],2'b0})+$signed({in[91],1'b0})+$signed({in[92],1'b0})+$signed(in[92])+$signed(-{in[118],3'b0})+$signed(-{in[119],3'b0})+$signed({in[63],1'b0})+$signed(sharing14_r)+$signed(-1);
assign weighted_sum[355] = $signed(-{in[120],3'b0})+$signed(-{in[121],3'b0})+$signed({in[65],1'b0})+$signed({in[66],2'b0})+$signed(-{in[122],1'b0})+$signed(in[66])+$signed(-{in[92],2'b0})+$signed({in[93],1'b0})+$signed({in[94],1'b0})+$signed(in[94])+$signed(sharing15_r)+$signed(-1);
assign weighted_sum[356] = $signed({in[96],1'b0})+$signed(in[96])+$signed(-{in[122],3'b0})+$signed(-{in[123],3'b0})+$signed({in[67],1'b0})+$signed({in[68],2'b0})+$signed(-{in[124],1'b0})+$signed(in[68])+$signed(-{in[94],2'b0})+$signed({in[95],1'b0})+$signed(sharing16_r)+$signed(-1);
assign weighted_sum[357] = $signed(-{in[96],2'b0})+$signed({in[97],1'b0})+$signed({in[98],1'b0})+$signed(in[98])+$signed(-{in[124],3'b0})+$signed(-{in[125],3'b0})+$signed({in[69],1'b0})+$signed({in[70],2'b0})+$signed(-{in[126],1'b0})+$signed(in[70])+$signed(sharing17_r)+$signed(-1);
assign weighted_sum[358] = $signed({in[72],2'b0})+$signed(-{in[128],1'b0})+$signed(in[72])+$signed(-{in[98],2'b0})+$signed({in[99],1'b0})+$signed({in[100],1'b0})+$signed(in[100])+$signed(-{in[126],3'b0})+$signed(-{in[127],3'b0})+$signed({in[71],1'b0})+$signed(sharing18_r)+$signed(-1);
assign weighted_sum[359] = $signed(-{in[128],3'b0})+$signed(-{in[129],3'b0})+$signed({in[73],1'b0})+$signed({in[74],2'b0})+$signed(-{in[130],1'b0})+$signed(in[74])+$signed(-{in[100],2'b0})+$signed({in[101],1'b0})+$signed({in[102],1'b0})+$signed(in[102])+$signed(sharing19_r)+$signed(-1);
assign weighted_sum[360] = $signed({in[104],1'b0})+$signed(in[104])+$signed(-{in[130],3'b0})+$signed(-{in[131],3'b0})+$signed({in[75],1'b0})+$signed({in[76],2'b0})+$signed(-{in[132],1'b0})+$signed(in[76])+$signed(-{in[102],2'b0})+$signed({in[103],1'b0})+$signed(sharing150_r)+$signed(-1);
assign weighted_sum[361] = $signed(-{in[104],2'b0})+$signed({in[105],1'b0})+$signed({in[106],1'b0})+$signed(in[106])+$signed(-{in[132],3'b0})+$signed(-{in[133],3'b0})+$signed({in[77],1'b0})+$signed({in[78],2'b0})+$signed(-{in[134],1'b0})+$signed(in[78])+$signed(sharing20_r)+$signed(-1);
assign weighted_sum[362] = $signed({in[80],2'b0})+$signed(-{in[136],1'b0})+$signed(in[80])+$signed(-{in[106],2'b0})+$signed({in[107],1'b0})+$signed({in[108],1'b0})+$signed(in[108])+$signed(-{in[134],3'b0})+$signed(-{in[135],3'b0})+$signed({in[79],1'b0})+$signed(sharing21_r)+$signed(-1);
assign weighted_sum[363] = $signed(-{in[136],3'b0})+$signed(-{in[137],3'b0})+$signed({in[81],1'b0})+$signed({in[82],2'b0})+$signed(-{in[138],1'b0})+$signed(in[82])+$signed(-{in[108],2'b0})+$signed({in[109],1'b0})+$signed({in[110],1'b0})+$signed(in[110])+$signed(sharing22_r)+$signed(-1);
assign weighted_sum[364] = $signed(-{in[168],3'b0})+$signed(-{in[169],3'b0})+$signed({in[113],1'b0})+$signed({in[114],2'b0})+$signed(-{in[170],1'b0})+$signed(in[114])+$signed(-{in[140],2'b0})+$signed({in[141],1'b0})+$signed({in[142],1'b0})+$signed(in[142])+$signed(sharing23_r)+$signed(-1);
assign weighted_sum[365] = $signed({in[144],1'b0})+$signed(in[144])+$signed(-{in[170],3'b0})+$signed(-{in[171],3'b0})+$signed({in[115],1'b0})+$signed({in[116],2'b0})+$signed(-{in[172],1'b0})+$signed(in[116])+$signed(-{in[142],2'b0})+$signed({in[143],1'b0})+$signed(sharing24_r)+$signed(-1);
assign weighted_sum[366] = $signed(-{in[144],2'b0})+$signed({in[145],1'b0})+$signed({in[146],1'b0})+$signed(in[146])+$signed(-{in[172],3'b0})+$signed(-{in[173],3'b0})+$signed({in[117],1'b0})+$signed({in[118],2'b0})+$signed(-{in[174],1'b0})+$signed(in[118])+$signed(sharing25_r)+$signed(-1);
assign weighted_sum[367] = $signed({in[120],2'b0})+$signed(-{in[176],1'b0})+$signed(in[120])+$signed(-{in[146],2'b0})+$signed({in[147],1'b0})+$signed({in[148],1'b0})+$signed(in[148])+$signed(-{in[174],3'b0})+$signed(-{in[175],3'b0})+$signed({in[119],1'b0})+$signed(sharing26_r)+$signed(-1);
assign weighted_sum[368] = $signed(-{in[176],3'b0})+$signed(-{in[177],3'b0})+$signed({in[121],1'b0})+$signed({in[122],2'b0})+$signed(-{in[178],1'b0})+$signed(in[122])+$signed(-{in[148],2'b0})+$signed({in[149],1'b0})+$signed({in[150],1'b0})+$signed(in[150])+$signed(sharing151_r)+$signed(-1);
assign weighted_sum[369] = $signed({in[152],1'b0})+$signed(in[152])+$signed(-{in[178],3'b0})+$signed(-{in[179],3'b0})+$signed({in[123],1'b0})+$signed({in[124],2'b0})+$signed(-{in[180],1'b0})+$signed(in[124])+$signed(-{in[150],2'b0})+$signed({in[151],1'b0})+$signed(sharing27_r)+$signed(-1);
assign weighted_sum[370] = $signed(-{in[152],2'b0})+$signed({in[153],1'b0})+$signed({in[154],1'b0})+$signed(in[154])+$signed(-{in[180],3'b0})+$signed(-{in[181],3'b0})+$signed({in[125],1'b0})+$signed({in[126],2'b0})+$signed(-{in[182],1'b0})+$signed(in[126])+$signed(sharing28_r)+$signed(-1);
assign weighted_sum[371] = $signed({in[128],2'b0})+$signed(-{in[184],1'b0})+$signed(in[128])+$signed(-{in[154],2'b0})+$signed({in[155],1'b0})+$signed({in[156],1'b0})+$signed(in[156])+$signed(-{in[182],3'b0})+$signed(-{in[183],3'b0})+$signed({in[127],1'b0})+$signed(sharing29_r)+$signed(-1);
assign weighted_sum[372] = $signed(-{in[184],3'b0})+$signed(-{in[185],3'b0})+$signed({in[129],1'b0})+$signed({in[130],2'b0})+$signed(-{in[186],1'b0})+$signed(in[130])+$signed(-{in[156],2'b0})+$signed({in[157],1'b0})+$signed({in[158],1'b0})+$signed(in[158])+$signed(sharing30_r)+$signed(-1);
assign weighted_sum[373] = $signed({in[160],1'b0})+$signed(in[160])+$signed(-{in[186],3'b0})+$signed(-{in[187],3'b0})+$signed({in[131],1'b0})+$signed({in[132],2'b0})+$signed(-{in[188],1'b0})+$signed(in[132])+$signed(-{in[158],2'b0})+$signed({in[159],1'b0})+$signed(sharing31_r)+$signed(-1);
assign weighted_sum[374] = $signed(-{in[160],2'b0})+$signed({in[161],1'b0})+$signed({in[162],1'b0})+$signed(in[162])+$signed(-{in[188],3'b0})+$signed(-{in[189],3'b0})+$signed({in[133],1'b0})+$signed({in[134],2'b0})+$signed(-{in[190],1'b0})+$signed(in[134])+$signed(sharing32_r)+$signed(-1);
assign weighted_sum[375] = $signed({in[136],2'b0})+$signed(-{in[192],1'b0})+$signed(in[136])+$signed(-{in[162],2'b0})+$signed({in[163],1'b0})+$signed({in[164],1'b0})+$signed(in[164])+$signed(-{in[190],3'b0})+$signed(-{in[191],3'b0})+$signed({in[135],1'b0})+$signed(sharing33_r)+$signed(-1);
assign weighted_sum[376] = $signed(-{in[192],3'b0})+$signed(-{in[193],3'b0})+$signed({in[137],1'b0})+$signed({in[138],2'b0})+$signed(-{in[194],1'b0})+$signed(in[138])+$signed(-{in[164],2'b0})+$signed({in[165],1'b0})+$signed({in[166],1'b0})+$signed(in[166])+$signed(sharing152_r)+$signed(-1);
assign weighted_sum[377] = $signed(-{in[224],3'b0})+$signed(-{in[225],3'b0})+$signed({in[169],1'b0})+$signed({in[170],2'b0})+$signed(-{in[226],1'b0})+$signed(in[170])+$signed(-{in[196],2'b0})+$signed({in[197],1'b0})+$signed({in[198],1'b0})+$signed(in[198])+$signed(sharing34_r)+$signed(-1);
assign weighted_sum[378] = $signed({in[200],1'b0})+$signed(in[200])+$signed(-{in[226],3'b0})+$signed(-{in[227],3'b0})+$signed({in[171],1'b0})+$signed({in[172],2'b0})+$signed(-{in[228],1'b0})+$signed(in[172])+$signed(-{in[198],2'b0})+$signed({in[199],1'b0})+$signed(sharing35_r)+$signed(-1);
assign weighted_sum[379] = $signed(-{in[200],2'b0})+$signed({in[201],1'b0})+$signed({in[202],1'b0})+$signed(in[202])+$signed(-{in[228],3'b0})+$signed(-{in[229],3'b0})+$signed({in[173],1'b0})+$signed({in[174],2'b0})+$signed(-{in[230],1'b0})+$signed(in[174])+$signed(sharing36_r)+$signed(-1);
assign weighted_sum[380] = $signed({in[176],2'b0})+$signed(-{in[232],1'b0})+$signed(in[176])+$signed(-{in[202],2'b0})+$signed({in[203],1'b0})+$signed({in[204],1'b0})+$signed(in[204])+$signed(-{in[230],3'b0})+$signed(-{in[231],3'b0})+$signed({in[175],1'b0})+$signed(sharing37_r)+$signed(-1);
assign weighted_sum[381] = $signed(-{in[232],3'b0})+$signed(-{in[233],3'b0})+$signed({in[177],1'b0})+$signed({in[178],2'b0})+$signed(-{in[234],1'b0})+$signed(in[178])+$signed(-{in[204],2'b0})+$signed({in[205],1'b0})+$signed({in[206],1'b0})+$signed(in[206])+$signed(sharing38_r)+$signed(-1);
assign weighted_sum[382] = $signed({in[208],1'b0})+$signed(in[208])+$signed(-{in[234],3'b0})+$signed(-{in[235],3'b0})+$signed({in[179],1'b0})+$signed({in[180],2'b0})+$signed(-{in[236],1'b0})+$signed(in[180])+$signed(-{in[206],2'b0})+$signed({in[207],1'b0})+$signed(sharing39_r)+$signed(-1);
assign weighted_sum[383] = $signed(-{in[208],2'b0})+$signed({in[209],1'b0})+$signed({in[210],1'b0})+$signed(in[210])+$signed(-{in[236],3'b0})+$signed(-{in[237],3'b0})+$signed({in[181],1'b0})+$signed({in[182],2'b0})+$signed(-{in[238],1'b0})+$signed(in[182])+$signed(sharing40_r)+$signed(-1);
assign weighted_sum[384] = $signed({in[184],2'b0})+$signed(-{in[240],1'b0})+$signed(in[184])+$signed(-{in[210],2'b0})+$signed({in[211],1'b0})+$signed({in[212],1'b0})+$signed(in[212])+$signed(-{in[238],3'b0})+$signed(-{in[239],3'b0})+$signed({in[183],1'b0})+$signed(sharing153_r)+$signed(-1);
assign weighted_sum[385] = $signed(-{in[240],3'b0})+$signed(-{in[241],3'b0})+$signed({in[185],1'b0})+$signed({in[186],2'b0})+$signed(-{in[242],1'b0})+$signed(in[186])+$signed(-{in[212],2'b0})+$signed({in[213],1'b0})+$signed({in[214],1'b0})+$signed(in[214])+$signed(sharing41_r)+$signed(-1);
assign weighted_sum[386] = $signed({in[216],1'b0})+$signed(in[216])+$signed(-{in[242],3'b0})+$signed(-{in[243],3'b0})+$signed({in[187],1'b0})+$signed({in[188],2'b0})+$signed(-{in[244],1'b0})+$signed(in[188])+$signed(-{in[214],2'b0})+$signed({in[215],1'b0})+$signed(sharing42_r)+$signed(-1);
assign weighted_sum[387] = $signed(-{in[216],2'b0})+$signed({in[217],1'b0})+$signed({in[218],1'b0})+$signed(in[218])+$signed(-{in[244],3'b0})+$signed(-{in[245],3'b0})+$signed({in[189],1'b0})+$signed({in[190],2'b0})+$signed(-{in[246],1'b0})+$signed(in[190])+$signed(sharing43_r)+$signed(-1);
assign weighted_sum[388] = $signed({in[192],2'b0})+$signed(-{in[248],1'b0})+$signed(in[192])+$signed(-{in[218],2'b0})+$signed({in[219],1'b0})+$signed({in[220],1'b0})+$signed(in[220])+$signed(-{in[246],3'b0})+$signed(-{in[247],3'b0})+$signed({in[191],1'b0})+$signed(sharing44_r)+$signed(-1);
assign weighted_sum[389] = $signed(-{in[248],3'b0})+$signed(-{in[249],3'b0})+$signed({in[193],1'b0})+$signed({in[194],2'b0})+$signed(-{in[250],1'b0})+$signed(in[194])+$signed(-{in[220],2'b0})+$signed({in[221],1'b0})+$signed({in[222],1'b0})+$signed(in[222])+$signed(sharing45_r)+$signed(-1);
assign weighted_sum[390] = $signed(-{in[280],3'b0})+$signed(-{in[281],3'b0})+$signed({in[225],1'b0})+$signed({in[226],2'b0})+$signed(-{in[282],1'b0})+$signed(in[226])+$signed(-{in[252],2'b0})+$signed({in[253],1'b0})+$signed({in[254],1'b0})+$signed(in[254])+$signed(sharing46_r)+$signed(-1);
assign weighted_sum[391] = $signed({in[256],1'b0})+$signed(in[256])+$signed(-{in[282],3'b0})+$signed(-{in[283],3'b0})+$signed({in[227],1'b0})+$signed({in[228],2'b0})+$signed(-{in[284],1'b0})+$signed(in[228])+$signed(-{in[254],2'b0})+$signed({in[255],1'b0})+$signed(sharing47_r)+$signed(-1);
assign weighted_sum[392] = $signed(-{in[256],2'b0})+$signed({in[257],1'b0})+$signed({in[258],1'b0})+$signed(in[258])+$signed(-{in[284],3'b0})+$signed(-{in[285],3'b0})+$signed({in[229],1'b0})+$signed({in[230],2'b0})+$signed(-{in[286],1'b0})+$signed(in[230])+$signed(sharing154_r)+$signed(-1);
assign weighted_sum[393] = $signed({in[232],2'b0})+$signed(-{in[288],1'b0})+$signed(in[232])+$signed(-{in[258],2'b0})+$signed({in[259],1'b0})+$signed({in[260],1'b0})+$signed(in[260])+$signed(-{in[286],3'b0})+$signed(-{in[287],3'b0})+$signed({in[231],1'b0})+$signed(sharing48_r)+$signed(-1);
assign weighted_sum[394] = $signed(-{in[288],3'b0})+$signed(-{in[289],3'b0})+$signed({in[233],1'b0})+$signed({in[234],2'b0})+$signed(-{in[290],1'b0})+$signed(in[234])+$signed(-{in[260],2'b0})+$signed({in[261],1'b0})+$signed({in[262],1'b0})+$signed(in[262])+$signed(sharing49_r)+$signed(-1);
assign weighted_sum[395] = $signed({in[264],1'b0})+$signed(in[264])+$signed(-{in[290],3'b0})+$signed(-{in[291],3'b0})+$signed({in[235],1'b0})+$signed({in[236],2'b0})+$signed(-{in[292],1'b0})+$signed(in[236])+$signed(-{in[262],2'b0})+$signed({in[263],1'b0})+$signed(sharing50_r)+$signed(-1);
assign weighted_sum[396] = $signed(-{in[264],2'b0})+$signed({in[265],1'b0})+$signed({in[266],1'b0})+$signed(in[266])+$signed(-{in[292],3'b0})+$signed(-{in[293],3'b0})+$signed({in[237],1'b0})+$signed({in[238],2'b0})+$signed(-{in[294],1'b0})+$signed(in[238])+$signed(sharing51_r)+$signed(-1);
assign weighted_sum[397] = $signed({in[240],2'b0})+$signed(-{in[296],1'b0})+$signed(in[240])+$signed(-{in[266],2'b0})+$signed({in[267],1'b0})+$signed({in[268],1'b0})+$signed(in[268])+$signed(-{in[294],3'b0})+$signed(-{in[295],3'b0})+$signed({in[239],1'b0})+$signed(sharing52_r)+$signed(-1);
assign weighted_sum[398] = $signed(-{in[296],3'b0})+$signed(-{in[297],3'b0})+$signed({in[241],1'b0})+$signed({in[242],2'b0})+$signed(-{in[298],1'b0})+$signed(in[242])+$signed(-{in[268],2'b0})+$signed({in[269],1'b0})+$signed({in[270],1'b0})+$signed(in[270])+$signed(sharing53_r)+$signed(-1);
assign weighted_sum[399] = $signed({in[272],1'b0})+$signed(in[272])+$signed(-{in[298],3'b0})+$signed(-{in[299],3'b0})+$signed({in[243],1'b0})+$signed({in[244],2'b0})+$signed(-{in[300],1'b0})+$signed(in[244])+$signed(-{in[270],2'b0})+$signed({in[271],1'b0})+$signed(sharing54_r)+$signed(-1);
assign weighted_sum[400] = $signed(-{in[272],2'b0})+$signed({in[273],1'b0})+$signed({in[274],1'b0})+$signed(in[274])+$signed(-{in[300],3'b0})+$signed(-{in[301],3'b0})+$signed({in[245],1'b0})+$signed({in[246],2'b0})+$signed(-{in[302],1'b0})+$signed(in[246])+$signed(sharing155_r)+$signed(-1);
assign weighted_sum[401] = $signed({in[248],2'b0})+$signed(-{in[304],1'b0})+$signed(in[248])+$signed(-{in[274],2'b0})+$signed({in[275],1'b0})+$signed({in[276],1'b0})+$signed(in[276])+$signed(-{in[302],3'b0})+$signed(-{in[303],3'b0})+$signed({in[247],1'b0})+$signed(sharing55_r)+$signed(-1);
assign weighted_sum[402] = $signed(-{in[304],3'b0})+$signed(-{in[305],3'b0})+$signed({in[249],1'b0})+$signed({in[250],2'b0})+$signed(-{in[306],1'b0})+$signed(in[250])+$signed(-{in[276],2'b0})+$signed({in[277],1'b0})+$signed({in[278],1'b0})+$signed(in[278])+$signed(sharing56_r)+$signed(-1);
assign weighted_sum[403] = $signed(-{in[336],3'b0})+$signed(-{in[337],3'b0})+$signed({in[281],1'b0})+$signed({in[282],2'b0})+$signed(-{in[338],1'b0})+$signed(in[282])+$signed(-{in[308],2'b0})+$signed({in[309],1'b0})+$signed({in[310],1'b0})+$signed(in[310])+$signed(sharing57_r)+$signed(-1);
assign weighted_sum[404] = $signed({in[312],1'b0})+$signed(in[312])+$signed(-{in[338],3'b0})+$signed(-{in[339],3'b0})+$signed({in[283],1'b0})+$signed({in[284],2'b0})+$signed(-{in[340],1'b0})+$signed(in[284])+$signed(-{in[310],2'b0})+$signed({in[311],1'b0})+$signed(sharing58_r)+$signed(-1);
assign weighted_sum[405] = $signed(-{in[312],2'b0})+$signed({in[313],1'b0})+$signed({in[314],1'b0})+$signed(in[314])+$signed(-{in[340],3'b0})+$signed(-{in[341],3'b0})+$signed({in[285],1'b0})+$signed({in[286],2'b0})+$signed(-{in[342],1'b0})+$signed(in[286])+$signed(sharing59_r)+$signed(-1);
assign weighted_sum[406] = $signed({in[288],2'b0})+$signed(-{in[344],1'b0})+$signed(in[288])+$signed(-{in[314],2'b0})+$signed({in[315],1'b0})+$signed({in[316],1'b0})+$signed(in[316])+$signed(-{in[342],3'b0})+$signed(-{in[343],3'b0})+$signed({in[287],1'b0})+$signed(sharing60_r)+$signed(-1);
assign weighted_sum[407] = $signed(-{in[344],3'b0})+$signed(-{in[345],3'b0})+$signed({in[289],1'b0})+$signed({in[290],2'b0})+$signed(-{in[346],1'b0})+$signed(in[290])+$signed(-{in[316],2'b0})+$signed({in[317],1'b0})+$signed({in[318],1'b0})+$signed(in[318])+$signed(sharing61_r)+$signed(-1);
assign weighted_sum[408] = $signed({in[320],1'b0})+$signed(in[320])+$signed(-{in[346],3'b0})+$signed(-{in[347],3'b0})+$signed({in[291],1'b0})+$signed({in[292],2'b0})+$signed(-{in[348],1'b0})+$signed(in[292])+$signed(-{in[318],2'b0})+$signed({in[319],1'b0})+$signed(sharing156_r)+$signed(-1);
assign weighted_sum[409] = $signed(-{in[320],2'b0})+$signed({in[321],1'b0})+$signed({in[322],1'b0})+$signed(in[322])+$signed(-{in[348],3'b0})+$signed(-{in[349],3'b0})+$signed({in[293],1'b0})+$signed({in[294],2'b0})+$signed(-{in[350],1'b0})+$signed(in[294])+$signed(sharing62_r)+$signed(-1);
assign weighted_sum[410] = $signed({in[296],2'b0})+$signed(-{in[352],1'b0})+$signed(in[296])+$signed(-{in[322],2'b0})+$signed({in[323],1'b0})+$signed({in[324],1'b0})+$signed(in[324])+$signed(-{in[350],3'b0})+$signed(-{in[351],3'b0})+$signed({in[295],1'b0})+$signed(sharing63_r)+$signed(-1);
assign weighted_sum[411] = $signed(-{in[352],3'b0})+$signed(-{in[353],3'b0})+$signed({in[297],1'b0})+$signed({in[298],2'b0})+$signed(-{in[354],1'b0})+$signed(in[298])+$signed(-{in[324],2'b0})+$signed({in[325],1'b0})+$signed({in[326],1'b0})+$signed(in[326])+$signed(sharing64_r)+$signed(-1);
assign weighted_sum[412] = $signed({in[328],1'b0})+$signed(in[328])+$signed(-{in[354],3'b0})+$signed(-{in[355],3'b0})+$signed({in[299],1'b0})+$signed({in[300],2'b0})+$signed(-{in[356],1'b0})+$signed(in[300])+$signed(-{in[326],2'b0})+$signed({in[327],1'b0})+$signed(sharing65_r)+$signed(-1);
assign weighted_sum[413] = $signed(-{in[328],2'b0})+$signed({in[329],1'b0})+$signed({in[330],1'b0})+$signed(in[330])+$signed(-{in[356],3'b0})+$signed(-{in[357],3'b0})+$signed({in[301],1'b0})+$signed({in[302],2'b0})+$signed(-{in[358],1'b0})+$signed(in[302])+$signed(sharing66_r)+$signed(-1);
assign weighted_sum[414] = $signed({in[304],2'b0})+$signed(-{in[360],1'b0})+$signed(in[304])+$signed(-{in[330],2'b0})+$signed({in[331],1'b0})+$signed({in[332],1'b0})+$signed(in[332])+$signed(-{in[358],3'b0})+$signed(-{in[359],3'b0})+$signed({in[303],1'b0})+$signed(sharing67_r)+$signed(-1);
assign weighted_sum[415] = $signed(-{in[360],3'b0})+$signed(-{in[361],3'b0})+$signed({in[305],1'b0})+$signed({in[306],2'b0})+$signed(-{in[362],1'b0})+$signed(in[306])+$signed(-{in[332],2'b0})+$signed({in[333],1'b0})+$signed({in[334],1'b0})+$signed(in[334])+$signed(sharing68_r)+$signed(-1);
assign weighted_sum[416] = $signed(-{in[392],3'b0})+$signed(-{in[393],3'b0})+$signed({in[337],1'b0})+$signed({in[338],2'b0})+$signed(-{in[394],1'b0})+$signed(in[338])+$signed(-{in[364],2'b0})+$signed({in[365],1'b0})+$signed({in[366],1'b0})+$signed(in[366])+$signed(sharing157_r)+$signed(-1);
assign weighted_sum[417] = $signed({in[368],1'b0})+$signed(in[368])+$signed(-{in[394],3'b0})+$signed(-{in[395],3'b0})+$signed({in[339],1'b0})+$signed({in[340],2'b0})+$signed(-{in[396],1'b0})+$signed(in[340])+$signed(-{in[366],2'b0})+$signed({in[367],1'b0})+$signed(sharing69_r)+$signed(-1);
assign weighted_sum[418] = $signed(-{in[368],2'b0})+$signed({in[369],1'b0})+$signed({in[370],1'b0})+$signed(in[370])+$signed(-{in[396],3'b0})+$signed(-{in[397],3'b0})+$signed({in[341],1'b0})+$signed({in[342],2'b0})+$signed(-{in[398],1'b0})+$signed(in[342])+$signed(sharing70_r)+$signed(-1);
assign weighted_sum[419] = $signed({in[344],2'b0})+$signed(-{in[400],1'b0})+$signed(in[344])+$signed(-{in[370],2'b0})+$signed({in[371],1'b0})+$signed({in[372],1'b0})+$signed(in[372])+$signed(-{in[398],3'b0})+$signed(-{in[399],3'b0})+$signed({in[343],1'b0})+$signed(sharing71_r)+$signed(-1);
assign weighted_sum[420] = $signed(-{in[400],3'b0})+$signed(-{in[401],3'b0})+$signed({in[345],1'b0})+$signed({in[346],2'b0})+$signed(-{in[402],1'b0})+$signed(in[346])+$signed(-{in[372],2'b0})+$signed({in[373],1'b0})+$signed({in[374],1'b0})+$signed(in[374])+$signed(sharing72_r)+$signed(-1);
assign weighted_sum[421] = $signed({in[376],1'b0})+$signed(in[376])+$signed(-{in[402],3'b0})+$signed(-{in[403],3'b0})+$signed({in[347],1'b0})+$signed({in[348],2'b0})+$signed(-{in[404],1'b0})+$signed(in[348])+$signed(-{in[374],2'b0})+$signed({in[375],1'b0})+$signed(sharing73_r)+$signed(-1);
assign weighted_sum[422] = $signed(-{in[376],2'b0})+$signed({in[377],1'b0})+$signed({in[378],1'b0})+$signed(in[378])+$signed(-{in[404],3'b0})+$signed(-{in[405],3'b0})+$signed({in[349],1'b0})+$signed({in[350],2'b0})+$signed(-{in[406],1'b0})+$signed(in[350])+$signed(sharing74_r)+$signed(-1);
assign weighted_sum[423] = $signed({in[352],2'b0})+$signed(-{in[408],1'b0})+$signed(in[352])+$signed(-{in[378],2'b0})+$signed({in[379],1'b0})+$signed({in[380],1'b0})+$signed(in[380])+$signed(-{in[406],3'b0})+$signed(-{in[407],3'b0})+$signed({in[351],1'b0})+$signed(sharing75_r)+$signed(-1);
assign weighted_sum[424] = $signed(-{in[408],3'b0})+$signed(-{in[409],3'b0})+$signed({in[353],1'b0})+$signed({in[354],2'b0})+$signed(-{in[410],1'b0})+$signed(in[354])+$signed(-{in[380],2'b0})+$signed({in[381],1'b0})+$signed({in[382],1'b0})+$signed(in[382])+$signed(sharing158_r)+$signed(-1);
assign weighted_sum[425] = $signed({in[384],1'b0})+$signed(in[384])+$signed(-{in[410],3'b0})+$signed(-{in[411],3'b0})+$signed({in[355],1'b0})+$signed({in[356],2'b0})+$signed(-{in[412],1'b0})+$signed(in[356])+$signed(-{in[382],2'b0})+$signed({in[383],1'b0})+$signed(sharing76_r)+$signed(-1);
assign weighted_sum[426] = $signed(-{in[384],2'b0})+$signed({in[385],1'b0})+$signed({in[386],1'b0})+$signed(in[386])+$signed(-{in[412],3'b0})+$signed(-{in[413],3'b0})+$signed({in[357],1'b0})+$signed({in[358],2'b0})+$signed(-{in[414],1'b0})+$signed(in[358])+$signed(sharing77_r)+$signed(-1);
assign weighted_sum[427] = $signed({in[360],2'b0})+$signed(-{in[416],1'b0})+$signed(in[360])+$signed(-{in[386],2'b0})+$signed({in[387],1'b0})+$signed({in[388],1'b0})+$signed(in[388])+$signed(-{in[414],3'b0})+$signed(-{in[415],3'b0})+$signed({in[359],1'b0})+$signed(sharing78_r)+$signed(-1);
assign weighted_sum[428] = $signed(-{in[416],3'b0})+$signed(-{in[417],3'b0})+$signed({in[361],1'b0})+$signed({in[362],2'b0})+$signed(-{in[418],1'b0})+$signed(in[362])+$signed(-{in[388],2'b0})+$signed({in[389],1'b0})+$signed({in[390],1'b0})+$signed(in[390])+$signed(sharing79_r)+$signed(-1);
assign weighted_sum[429] = $signed(-{in[448],3'b0})+$signed(-{in[449],3'b0})+$signed({in[393],1'b0})+$signed({in[394],2'b0})+$signed(-{in[450],1'b0})+$signed(in[394])+$signed(-{in[420],2'b0})+$signed({in[421],1'b0})+$signed({in[422],1'b0})+$signed(in[422])+$signed(sharing80_r)+$signed(-1);
assign weighted_sum[430] = $signed({in[424],1'b0})+$signed(in[424])+$signed(-{in[450],3'b0})+$signed(-{in[451],3'b0})+$signed({in[395],1'b0})+$signed({in[396],2'b0})+$signed(-{in[452],1'b0})+$signed(in[396])+$signed(-{in[422],2'b0})+$signed({in[423],1'b0})+$signed(sharing81_r)+$signed(-1);
assign weighted_sum[431] = $signed(-{in[424],2'b0})+$signed({in[425],1'b0})+$signed({in[426],1'b0})+$signed(in[426])+$signed(-{in[452],3'b0})+$signed(-{in[453],3'b0})+$signed({in[397],1'b0})+$signed({in[398],2'b0})+$signed(-{in[454],1'b0})+$signed(in[398])+$signed(sharing82_r)+$signed(-1);
assign weighted_sum[432] = $signed({in[400],2'b0})+$signed(-{in[456],1'b0})+$signed(in[400])+$signed(-{in[426],2'b0})+$signed({in[427],1'b0})+$signed({in[428],1'b0})+$signed(in[428])+$signed(-{in[454],3'b0})+$signed(-{in[455],3'b0})+$signed({in[399],1'b0})+$signed(sharing159_r)+$signed(-1);
assign weighted_sum[433] = $signed(-{in[456],3'b0})+$signed(-{in[457],3'b0})+$signed({in[401],1'b0})+$signed({in[402],2'b0})+$signed(-{in[458],1'b0})+$signed(in[402])+$signed(-{in[428],2'b0})+$signed({in[429],1'b0})+$signed({in[430],1'b0})+$signed(in[430])+$signed(sharing83_r)+$signed(-1);
assign weighted_sum[434] = $signed({in[432],1'b0})+$signed(in[432])+$signed(-{in[458],3'b0})+$signed(-{in[459],3'b0})+$signed({in[403],1'b0})+$signed({in[404],2'b0})+$signed(-{in[460],1'b0})+$signed(in[404])+$signed(-{in[430],2'b0})+$signed({in[431],1'b0})+$signed(sharing84_r)+$signed(-1);
assign weighted_sum[435] = $signed(-{in[432],2'b0})+$signed({in[433],1'b0})+$signed({in[434],1'b0})+$signed(in[434])+$signed(-{in[460],3'b0})+$signed(-{in[461],3'b0})+$signed({in[405],1'b0})+$signed({in[406],2'b0})+$signed(-{in[462],1'b0})+$signed(in[406])+$signed(sharing85_r)+$signed(-1);
assign weighted_sum[436] = $signed({in[408],2'b0})+$signed(-{in[464],1'b0})+$signed(in[408])+$signed(-{in[434],2'b0})+$signed({in[435],1'b0})+$signed({in[436],1'b0})+$signed(in[436])+$signed(-{in[462],3'b0})+$signed(-{in[463],3'b0})+$signed({in[407],1'b0})+$signed(sharing86_r)+$signed(-1);
assign weighted_sum[437] = $signed(-{in[464],3'b0})+$signed(-{in[465],3'b0})+$signed({in[409],1'b0})+$signed({in[410],2'b0})+$signed(-{in[466],1'b0})+$signed(in[410])+$signed(-{in[436],2'b0})+$signed({in[437],1'b0})+$signed({in[438],1'b0})+$signed(in[438])+$signed(sharing87_r)+$signed(-1);
assign weighted_sum[438] = $signed({in[440],1'b0})+$signed(in[440])+$signed(-{in[466],3'b0})+$signed(-{in[467],3'b0})+$signed({in[411],1'b0})+$signed({in[412],2'b0})+$signed(-{in[468],1'b0})+$signed(in[412])+$signed(-{in[438],2'b0})+$signed({in[439],1'b0})+$signed(sharing88_r)+$signed(-1);
assign weighted_sum[439] = $signed(-{in[440],2'b0})+$signed({in[441],1'b0})+$signed({in[442],1'b0})+$signed(in[442])+$signed(-{in[468],3'b0})+$signed(-{in[469],3'b0})+$signed({in[413],1'b0})+$signed({in[414],2'b0})+$signed(-{in[470],1'b0})+$signed(in[414])+$signed(sharing89_r)+$signed(-1);
assign weighted_sum[440] = $signed({in[416],2'b0})+$signed(-{in[472],1'b0})+$signed(in[416])+$signed(-{in[442],2'b0})+$signed({in[443],1'b0})+$signed({in[444],1'b0})+$signed(in[444])+$signed(-{in[470],3'b0})+$signed(-{in[471],3'b0})+$signed({in[415],1'b0})+$signed(sharing160_r)+$signed(-1);
assign weighted_sum[441] = $signed(-{in[472],3'b0})+$signed(-{in[473],3'b0})+$signed({in[417],1'b0})+$signed({in[418],2'b0})+$signed(-{in[474],1'b0})+$signed(in[418])+$signed(-{in[444],2'b0})+$signed({in[445],1'b0})+$signed({in[446],1'b0})+$signed(in[446])+$signed(sharing90_r)+$signed(-1);
assign weighted_sum[442] = $signed(-{in[504],3'b0})+$signed(-{in[505],3'b0})+$signed({in[449],1'b0})+$signed({in[450],2'b0})+$signed(-{in[506],1'b0})+$signed(in[450])+$signed(-{in[476],2'b0})+$signed({in[477],1'b0})+$signed({in[478],1'b0})+$signed(in[478])+$signed(sharing91_r)+$signed(-1);
assign weighted_sum[443] = $signed({in[480],1'b0})+$signed(in[480])+$signed(-{in[506],3'b0})+$signed(-{in[507],3'b0})+$signed({in[451],1'b0})+$signed({in[452],2'b0})+$signed(-{in[508],1'b0})+$signed(in[452])+$signed(-{in[478],2'b0})+$signed({in[479],1'b0})+$signed(sharing92_r)+$signed(-1);
assign weighted_sum[444] = $signed(-{in[480],2'b0})+$signed({in[481],1'b0})+$signed({in[482],1'b0})+$signed(in[482])+$signed(-{in[508],3'b0})+$signed(-{in[509],3'b0})+$signed({in[453],1'b0})+$signed({in[454],2'b0})+$signed(-{in[510],1'b0})+$signed(in[454])+$signed(sharing93_r)+$signed(-1);
assign weighted_sum[445] = $signed({in[456],2'b0})+$signed(-{in[512],1'b0})+$signed(in[456])+$signed(-{in[482],2'b0})+$signed({in[483],1'b0})+$signed({in[484],1'b0})+$signed(in[484])+$signed(-{in[510],3'b0})+$signed(-{in[511],3'b0})+$signed({in[455],1'b0})+$signed(sharing94_r)+$signed(-1);
assign weighted_sum[446] = $signed(-{in[512],3'b0})+$signed(-{in[513],3'b0})+$signed({in[457],1'b0})+$signed({in[458],2'b0})+$signed(-{in[514],1'b0})+$signed(in[458])+$signed(-{in[484],2'b0})+$signed({in[485],1'b0})+$signed({in[486],1'b0})+$signed(in[486])+$signed(sharing95_r)+$signed(-1);
assign weighted_sum[447] = $signed({in[488],1'b0})+$signed(in[488])+$signed(-{in[514],3'b0})+$signed(-{in[515],3'b0})+$signed({in[459],1'b0})+$signed({in[460],2'b0})+$signed(-{in[516],1'b0})+$signed(in[460])+$signed(-{in[486],2'b0})+$signed({in[487],1'b0})+$signed(sharing96_r)+$signed(-1);
assign weighted_sum[448] = $signed(-{in[488],2'b0})+$signed({in[489],1'b0})+$signed({in[490],1'b0})+$signed(in[490])+$signed(-{in[516],3'b0})+$signed(-{in[517],3'b0})+$signed({in[461],1'b0})+$signed({in[462],2'b0})+$signed(-{in[518],1'b0})+$signed(in[462])+$signed(sharing161_r)+$signed(-1);
assign weighted_sum[449] = $signed({in[464],2'b0})+$signed(-{in[520],1'b0})+$signed(in[464])+$signed(-{in[490],2'b0})+$signed({in[491],1'b0})+$signed({in[492],1'b0})+$signed(in[492])+$signed(-{in[518],3'b0})+$signed(-{in[519],3'b0})+$signed({in[463],1'b0})+$signed(sharing97_r)+$signed(-1);
assign weighted_sum[450] = $signed(-{in[520],3'b0})+$signed(-{in[521],3'b0})+$signed({in[465],1'b0})+$signed({in[466],2'b0})+$signed(-{in[522],1'b0})+$signed(in[466])+$signed(-{in[492],2'b0})+$signed({in[493],1'b0})+$signed({in[494],1'b0})+$signed(in[494])+$signed(sharing98_r)+$signed(-1);
assign weighted_sum[451] = $signed({in[496],1'b0})+$signed(in[496])+$signed(-{in[522],3'b0})+$signed(-{in[523],3'b0})+$signed({in[467],1'b0})+$signed({in[468],2'b0})+$signed(-{in[524],1'b0})+$signed(in[468])+$signed(-{in[494],2'b0})+$signed({in[495],1'b0})+$signed(sharing99_r)+$signed(-1);
assign weighted_sum[452] = $signed(-{in[496],2'b0})+$signed({in[497],1'b0})+$signed({in[498],1'b0})+$signed(in[498])+$signed(-{in[524],3'b0})+$signed(-{in[525],3'b0})+$signed({in[469],1'b0})+$signed({in[470],2'b0})+$signed(-{in[526],1'b0})+$signed(in[470])+$signed(sharing100_r)+$signed(-1);
assign weighted_sum[453] = $signed({in[472],2'b0})+$signed(-{in[528],1'b0})+$signed(in[472])+$signed(-{in[498],2'b0})+$signed({in[499],1'b0})+$signed({in[500],1'b0})+$signed(in[500])+$signed(-{in[526],3'b0})+$signed(-{in[527],3'b0})+$signed({in[471],1'b0})+$signed(sharing101_r)+$signed(-1);
assign weighted_sum[454] = $signed(-{in[528],3'b0})+$signed(-{in[529],3'b0})+$signed({in[473],1'b0})+$signed({in[474],2'b0})+$signed(-{in[530],1'b0})+$signed(in[474])+$signed(-{in[500],2'b0})+$signed({in[501],1'b0})+$signed({in[502],1'b0})+$signed(in[502])+$signed(sharing102_r)+$signed(-1);
assign weighted_sum[455] = $signed(-{in[560],3'b0})+$signed(-{in[561],3'b0})+$signed({in[505],1'b0})+$signed({in[506],2'b0})+$signed(-{in[562],1'b0})+$signed(in[506])+$signed(-{in[532],2'b0})+$signed({in[533],1'b0})+$signed({in[534],1'b0})+$signed(in[534])+$signed(sharing103_r)+$signed(-1);
assign weighted_sum[456] = $signed({in[536],1'b0})+$signed(in[536])+$signed(-{in[562],3'b0})+$signed(-{in[563],3'b0})+$signed({in[507],1'b0})+$signed({in[508],2'b0})+$signed(-{in[564],1'b0})+$signed(in[508])+$signed(-{in[534],2'b0})+$signed({in[535],1'b0})+$signed(sharing162_r)+$signed(-1);
assign weighted_sum[457] = $signed(-{in[536],2'b0})+$signed({in[537],1'b0})+$signed({in[538],1'b0})+$signed(in[538])+$signed(-{in[564],3'b0})+$signed(-{in[565],3'b0})+$signed({in[509],1'b0})+$signed({in[510],2'b0})+$signed(-{in[566],1'b0})+$signed(in[510])+$signed(sharing104_r)+$signed(-1);
assign weighted_sum[458] = $signed({in[512],2'b0})+$signed(-{in[568],1'b0})+$signed(in[512])+$signed(-{in[538],2'b0})+$signed({in[539],1'b0})+$signed({in[540],1'b0})+$signed(in[540])+$signed(-{in[566],3'b0})+$signed(-{in[567],3'b0})+$signed({in[511],1'b0})+$signed(sharing105_r)+$signed(-1);
assign weighted_sum[459] = $signed(-{in[568],3'b0})+$signed(-{in[569],3'b0})+$signed({in[513],1'b0})+$signed({in[514],2'b0})+$signed(-{in[570],1'b0})+$signed(in[514])+$signed(-{in[540],2'b0})+$signed({in[541],1'b0})+$signed({in[542],1'b0})+$signed(in[542])+$signed(sharing106_r)+$signed(-1);
assign weighted_sum[460] = $signed({in[544],1'b0})+$signed(in[544])+$signed(-{in[570],3'b0})+$signed(-{in[571],3'b0})+$signed({in[515],1'b0})+$signed({in[516],2'b0})+$signed(-{in[572],1'b0})+$signed(in[516])+$signed(-{in[542],2'b0})+$signed({in[543],1'b0})+$signed(sharing107_r)+$signed(-1);
assign weighted_sum[461] = $signed(-{in[544],2'b0})+$signed({in[545],1'b0})+$signed({in[546],1'b0})+$signed(in[546])+$signed(-{in[572],3'b0})+$signed(-{in[573],3'b0})+$signed({in[517],1'b0})+$signed({in[518],2'b0})+$signed(-{in[574],1'b0})+$signed(in[518])+$signed(sharing108_r)+$signed(-1);
assign weighted_sum[462] = $signed({in[520],2'b0})+$signed(-{in[576],1'b0})+$signed(in[520])+$signed(-{in[546],2'b0})+$signed({in[547],1'b0})+$signed({in[548],1'b0})+$signed(in[548])+$signed(-{in[574],3'b0})+$signed(-{in[575],3'b0})+$signed({in[519],1'b0})+$signed(sharing109_r)+$signed(-1);
assign weighted_sum[463] = $signed(-{in[576],3'b0})+$signed(-{in[577],3'b0})+$signed({in[521],1'b0})+$signed({in[522],2'b0})+$signed(-{in[578],1'b0})+$signed(in[522])+$signed(-{in[548],2'b0})+$signed({in[549],1'b0})+$signed({in[550],1'b0})+$signed(in[550])+$signed(sharing110_r)+$signed(-1);
assign weighted_sum[464] = $signed({in[552],1'b0})+$signed(in[552])+$signed(-{in[578],3'b0})+$signed(-{in[579],3'b0})+$signed({in[523],1'b0})+$signed({in[524],2'b0})+$signed(-{in[580],1'b0})+$signed(in[524])+$signed(-{in[550],2'b0})+$signed({in[551],1'b0})+$signed(sharing163_r)+$signed(-1);
assign weighted_sum[465] = $signed(-{in[552],2'b0})+$signed({in[553],1'b0})+$signed({in[554],1'b0})+$signed(in[554])+$signed(-{in[580],3'b0})+$signed(-{in[581],3'b0})+$signed({in[525],1'b0})+$signed({in[526],2'b0})+$signed(-{in[582],1'b0})+$signed(in[526])+$signed(sharing111_r)+$signed(-1);
assign weighted_sum[466] = $signed({in[528],2'b0})+$signed(-{in[584],1'b0})+$signed(in[528])+$signed(-{in[554],2'b0})+$signed({in[555],1'b0})+$signed({in[556],1'b0})+$signed(in[556])+$signed(-{in[582],3'b0})+$signed(-{in[583],3'b0})+$signed({in[527],1'b0})+$signed(sharing112_r)+$signed(-1);
assign weighted_sum[467] = $signed(-{in[584],3'b0})+$signed(-{in[585],3'b0})+$signed({in[529],1'b0})+$signed({in[530],2'b0})+$signed(-{in[586],1'b0})+$signed(in[530])+$signed(-{in[556],2'b0})+$signed({in[557],1'b0})+$signed({in[558],1'b0})+$signed(in[558])+$signed(sharing113_r)+$signed(-1);
assign weighted_sum[468] = $signed(-{in[616],3'b0})+$signed(-{in[617],3'b0})+$signed({in[561],1'b0})+$signed({in[562],2'b0})+$signed(-{in[618],1'b0})+$signed(in[562])+$signed(-{in[588],2'b0})+$signed({in[589],1'b0})+$signed({in[590],1'b0})+$signed(in[590])+$signed(sharing114_r)+$signed(-1);
assign weighted_sum[469] = $signed({in[592],1'b0})+$signed(in[592])+$signed(-{in[618],3'b0})+$signed(-{in[619],3'b0})+$signed({in[563],1'b0})+$signed({in[564],2'b0})+$signed(-{in[620],1'b0})+$signed(in[564])+$signed(-{in[590],2'b0})+$signed({in[591],1'b0})+$signed(sharing115_r)+$signed(-1);
assign weighted_sum[470] = $signed(-{in[592],2'b0})+$signed({in[593],1'b0})+$signed({in[594],1'b0})+$signed(in[594])+$signed(-{in[620],3'b0})+$signed(-{in[621],3'b0})+$signed({in[565],1'b0})+$signed({in[566],2'b0})+$signed(-{in[622],1'b0})+$signed(in[566])+$signed(sharing116_r)+$signed(-1);
assign weighted_sum[471] = $signed({in[568],2'b0})+$signed(-{in[624],1'b0})+$signed(in[568])+$signed(-{in[594],2'b0})+$signed({in[595],1'b0})+$signed({in[596],1'b0})+$signed(in[596])+$signed(-{in[622],3'b0})+$signed(-{in[623],3'b0})+$signed({in[567],1'b0})+$signed(sharing117_r)+$signed(-1);
assign weighted_sum[472] = $signed(-{in[624],3'b0})+$signed(-{in[625],3'b0})+$signed({in[569],1'b0})+$signed({in[570],2'b0})+$signed(-{in[626],1'b0})+$signed(in[570])+$signed(-{in[596],2'b0})+$signed({in[597],1'b0})+$signed({in[598],1'b0})+$signed(in[598])+$signed(sharing164_r)+$signed(-1);
assign weighted_sum[473] = $signed({in[600],1'b0})+$signed(in[600])+$signed(-{in[626],3'b0})+$signed(-{in[627],3'b0})+$signed({in[571],1'b0})+$signed({in[572],2'b0})+$signed(-{in[628],1'b0})+$signed(in[572])+$signed(-{in[598],2'b0})+$signed({in[599],1'b0})+$signed(sharing118_r)+$signed(-1);
assign weighted_sum[474] = $signed(-{in[600],2'b0})+$signed({in[601],1'b0})+$signed({in[602],1'b0})+$signed(in[602])+$signed(-{in[628],3'b0})+$signed(-{in[629],3'b0})+$signed({in[573],1'b0})+$signed({in[574],2'b0})+$signed(-{in[630],1'b0})+$signed(in[574])+$signed(sharing119_r)+$signed(-1);
assign weighted_sum[475] = $signed({in[576],2'b0})+$signed(-{in[632],1'b0})+$signed(in[576])+$signed(-{in[602],2'b0})+$signed({in[603],1'b0})+$signed({in[604],1'b0})+$signed(in[604])+$signed(-{in[630],3'b0})+$signed(-{in[631],3'b0})+$signed({in[575],1'b0})+$signed(sharing120_r)+$signed(-1);
assign weighted_sum[476] = $signed(-{in[632],3'b0})+$signed(-{in[633],3'b0})+$signed({in[577],1'b0})+$signed({in[578],2'b0})+$signed(-{in[634],1'b0})+$signed(in[578])+$signed(-{in[604],2'b0})+$signed({in[605],1'b0})+$signed({in[606],1'b0})+$signed(in[606])+$signed(sharing121_r)+$signed(-1);
assign weighted_sum[477] = $signed({in[608],1'b0})+$signed(in[608])+$signed(-{in[634],3'b0})+$signed(-{in[635],3'b0})+$signed({in[579],1'b0})+$signed({in[580],2'b0})+$signed(-{in[636],1'b0})+$signed(in[580])+$signed(-{in[606],2'b0})+$signed({in[607],1'b0})+$signed(sharing122_r)+$signed(-1);
assign weighted_sum[478] = $signed(-{in[608],2'b0})+$signed({in[609],1'b0})+$signed({in[610],1'b0})+$signed(in[610])+$signed(-{in[636],3'b0})+$signed(-{in[637],3'b0})+$signed({in[581],1'b0})+$signed({in[582],2'b0})+$signed(-{in[638],1'b0})+$signed(in[582])+$signed(sharing123_r)+$signed(-1);
assign weighted_sum[479] = $signed({in[584],2'b0})+$signed(-{in[640],1'b0})+$signed(in[584])+$signed(-{in[610],2'b0})+$signed({in[611],1'b0})+$signed({in[612],1'b0})+$signed(in[612])+$signed(-{in[638],3'b0})+$signed(-{in[639],3'b0})+$signed({in[583],1'b0})+$signed(sharing124_r)+$signed(-1);
assign weighted_sum[480] = $signed(-{in[640],3'b0})+$signed(-{in[641],3'b0})+$signed({in[585],1'b0})+$signed({in[586],2'b0})+$signed(-{in[642],1'b0})+$signed(in[586])+$signed(-{in[612],2'b0})+$signed({in[613],1'b0})+$signed({in[614],1'b0})+$signed(in[614])+$signed(sharing165_r)+$signed(-1);
assign weighted_sum[481] = $signed(-{in[672],3'b0})+$signed(-{in[673],3'b0})+$signed({in[617],1'b0})+$signed({in[618],2'b0})+$signed(-{in[674],1'b0})+$signed(in[618])+$signed(-{in[644],2'b0})+$signed({in[645],1'b0})+$signed({in[646],1'b0})+$signed(in[646])+$signed(sharing125_r)+$signed(-1);
assign weighted_sum[482] = $signed({in[648],1'b0})+$signed(in[648])+$signed(-{in[674],3'b0})+$signed(-{in[675],3'b0})+$signed({in[619],1'b0})+$signed({in[620],2'b0})+$signed(-{in[676],1'b0})+$signed(in[620])+$signed(-{in[646],2'b0})+$signed({in[647],1'b0})+$signed(sharing126_r)+$signed(-1);
assign weighted_sum[483] = $signed(-{in[648],2'b0})+$signed({in[649],1'b0})+$signed({in[650],1'b0})+$signed(in[650])+$signed(-{in[676],3'b0})+$signed(-{in[677],3'b0})+$signed({in[621],1'b0})+$signed({in[622],2'b0})+$signed(-{in[678],1'b0})+$signed(in[622])+$signed(sharing127_r)+$signed(-1);
assign weighted_sum[484] = $signed({in[624],2'b0})+$signed(-{in[680],1'b0})+$signed(in[624])+$signed(-{in[650],2'b0})+$signed({in[651],1'b0})+$signed({in[652],1'b0})+$signed(in[652])+$signed(-{in[678],3'b0})+$signed(-{in[679],3'b0})+$signed({in[623],1'b0})+$signed(sharing128_r)+$signed(-1);
assign weighted_sum[485] = $signed(-{in[680],3'b0})+$signed(-{in[681],3'b0})+$signed({in[625],1'b0})+$signed({in[626],2'b0})+$signed(-{in[682],1'b0})+$signed(in[626])+$signed(-{in[652],2'b0})+$signed({in[653],1'b0})+$signed({in[654],1'b0})+$signed(in[654])+$signed(sharing129_r)+$signed(-1);
assign weighted_sum[486] = $signed({in[656],1'b0})+$signed(in[656])+$signed(-{in[682],3'b0})+$signed(-{in[683],3'b0})+$signed({in[627],1'b0})+$signed({in[628],2'b0})+$signed(-{in[684],1'b0})+$signed(in[628])+$signed(-{in[654],2'b0})+$signed({in[655],1'b0})+$signed(sharing130_r)+$signed(-1);
assign weighted_sum[487] = $signed(-{in[656],2'b0})+$signed({in[657],1'b0})+$signed({in[658],1'b0})+$signed(in[658])+$signed(-{in[684],3'b0})+$signed(-{in[685],3'b0})+$signed({in[629],1'b0})+$signed({in[630],2'b0})+$signed(-{in[686],1'b0})+$signed(in[630])+$signed(sharing131_r)+$signed(-1);
assign weighted_sum[488] = $signed({in[632],2'b0})+$signed(-{in[688],1'b0})+$signed(in[632])+$signed(-{in[658],2'b0})+$signed({in[659],1'b0})+$signed({in[660],1'b0})+$signed(in[660])+$signed(-{in[686],3'b0})+$signed(-{in[687],3'b0})+$signed({in[631],1'b0})+$signed(sharing166_r)+$signed(-1);
assign weighted_sum[489] = $signed(-{in[688],3'b0})+$signed(-{in[689],3'b0})+$signed({in[633],1'b0})+$signed({in[634],2'b0})+$signed(-{in[690],1'b0})+$signed(in[634])+$signed(-{in[660],2'b0})+$signed({in[661],1'b0})+$signed({in[662],1'b0})+$signed(in[662])+$signed(sharing132_r)+$signed(-1);
assign weighted_sum[490] = $signed({in[664],1'b0})+$signed(in[664])+$signed(-{in[690],3'b0})+$signed(-{in[691],3'b0})+$signed({in[635],1'b0})+$signed({in[636],2'b0})+$signed(-{in[692],1'b0})+$signed(in[636])+$signed(-{in[662],2'b0})+$signed({in[663],1'b0})+$signed(sharing133_r)+$signed(-1);
assign weighted_sum[491] = $signed(-{in[664],2'b0})+$signed({in[665],1'b0})+$signed({in[666],1'b0})+$signed(in[666])+$signed(-{in[692],3'b0})+$signed(-{in[693],3'b0})+$signed({in[637],1'b0})+$signed({in[638],2'b0})+$signed(-{in[694],1'b0})+$signed(in[638])+$signed(sharing134_r)+$signed(-1);
assign weighted_sum[492] = $signed({in[640],2'b0})+$signed(-{in[696],1'b0})+$signed(in[640])+$signed(-{in[666],2'b0})+$signed({in[667],1'b0})+$signed({in[668],1'b0})+$signed(in[668])+$signed(-{in[694],3'b0})+$signed(-{in[695],3'b0})+$signed({in[639],1'b0})+$signed(sharing135_r)+$signed(-1);
assign weighted_sum[493] = $signed(-{in[696],3'b0})+$signed(-{in[697],3'b0})+$signed({in[641],1'b0})+$signed({in[642],2'b0})+$signed(-{in[698],1'b0})+$signed(in[642])+$signed(-{in[668],2'b0})+$signed({in[669],1'b0})+$signed({in[670],1'b0})+$signed(in[670])+$signed(sharing136_r)+$signed(-1);
assign weighted_sum[494] = $signed(-{in[728],3'b0})+$signed(-{in[729],3'b0})+$signed({in[673],1'b0})+$signed({in[674],2'b0})+$signed(-{in[730],1'b0})+$signed(in[674])+$signed(-{in[700],2'b0})+$signed({in[701],1'b0})+$signed({in[702],1'b0})+$signed(in[702])+$signed(sharing137_r)+$signed(-1);
assign weighted_sum[495] = $signed({in[704],1'b0})+$signed(in[704])+$signed(-{in[730],3'b0})+$signed(-{in[731],3'b0})+$signed({in[675],1'b0})+$signed({in[676],2'b0})+$signed(-{in[732],1'b0})+$signed(in[676])+$signed(-{in[702],2'b0})+$signed({in[703],1'b0})+$signed(sharing138_r)+$signed(-1);
assign weighted_sum[496] = $signed(-{in[704],2'b0})+$signed({in[705],1'b0})+$signed({in[706],1'b0})+$signed(in[706])+$signed(-{in[732],3'b0})+$signed(-{in[733],3'b0})+$signed({in[677],1'b0})+$signed({in[678],2'b0})+$signed(-{in[734],1'b0})+$signed(in[678])+$signed(sharing167_r)+$signed(-1);
assign weighted_sum[497] = $signed({in[680],2'b0})+$signed(-{in[736],1'b0})+$signed(in[680])+$signed(-{in[706],2'b0})+$signed({in[707],1'b0})+$signed({in[708],1'b0})+$signed(in[708])+$signed(-{in[734],3'b0})+$signed(-{in[735],3'b0})+$signed({in[679],1'b0})+$signed(sharing139_r)+$signed(-1);
assign weighted_sum[498] = $signed(-{in[736],3'b0})+$signed(-{in[737],3'b0})+$signed({in[681],1'b0})+$signed({in[682],2'b0})+$signed(-{in[738],1'b0})+$signed(in[682])+$signed(-{in[708],2'b0})+$signed({in[709],1'b0})+$signed({in[710],1'b0})+$signed(in[710])+$signed(sharing140_r)+$signed(-1);
assign weighted_sum[499] = $signed({in[712],1'b0})+$signed(in[712])+$signed(-{in[738],3'b0})+$signed(-{in[739],3'b0})+$signed({in[683],1'b0})+$signed({in[684],2'b0})+$signed(-{in[740],1'b0})+$signed(in[684])+$signed(-{in[710],2'b0})+$signed({in[711],1'b0})+$signed(sharing141_r)+$signed(-1);
assign weighted_sum[500] = $signed(-{in[712],2'b0})+$signed({in[713],1'b0})+$signed({in[714],1'b0})+$signed(in[714])+$signed(-{in[740],3'b0})+$signed(-{in[741],3'b0})+$signed({in[685],1'b0})+$signed({in[686],2'b0})+$signed(-{in[742],1'b0})+$signed(in[686])+$signed(sharing142_r)+$signed(-1);
assign weighted_sum[501] = $signed({in[688],2'b0})+$signed(-{in[744],1'b0})+$signed(in[688])+$signed(-{in[714],2'b0})+$signed({in[715],1'b0})+$signed({in[716],1'b0})+$signed(in[716])+$signed(-{in[742],3'b0})+$signed(-{in[743],3'b0})+$signed({in[687],1'b0})+$signed(sharing143_r)+$signed(-1);
assign weighted_sum[502] = $signed(-{in[744],3'b0})+$signed(-{in[745],3'b0})+$signed({in[689],1'b0})+$signed({in[690],2'b0})+$signed(-{in[746],1'b0})+$signed(in[690])+$signed(-{in[716],2'b0})+$signed({in[717],1'b0})+$signed({in[718],1'b0})+$signed(in[718])+$signed(sharing144_r)+$signed(-1);
assign weighted_sum[503] = $signed({in[720],1'b0})+$signed(in[720])+$signed(-{in[746],3'b0})+$signed(-{in[747],3'b0})+$signed({in[691],1'b0})+$signed({in[692],2'b0})+$signed(-{in[748],1'b0})+$signed(in[692])+$signed(-{in[718],2'b0})+$signed({in[719],1'b0})+$signed(sharing145_r)+$signed(-1);
assign weighted_sum[504] = $signed(-{in[720],2'b0})+$signed({in[721],1'b0})+$signed({in[722],1'b0})+$signed(in[722])+$signed(-{in[748],3'b0})+$signed(-{in[749],3'b0})+$signed({in[693],1'b0})+$signed({in[694],2'b0})+$signed(-{in[750],1'b0})+$signed(in[694])+$signed(sharing168_r)+$signed(-1);
assign weighted_sum[505] = $signed({in[696],2'b0})+$signed(-{in[752],1'b0})+$signed(in[696])+$signed(-{in[722],2'b0})+$signed({in[723],1'b0})+$signed({in[724],1'b0})+$signed(in[724])+$signed(-{in[750],3'b0})+$signed(-{in[751],3'b0})+$signed({in[695],1'b0})+$signed(sharing146_r)+$signed(-1);
assign weighted_sum[506] = $signed(-{in[752],3'b0})+$signed(-{in[753],3'b0})+$signed({in[697],1'b0})+$signed({in[698],2'b0})+$signed(-{in[754],1'b0})+$signed(in[698])+$signed(-{in[724],2'b0})+$signed({in[725],1'b0})+$signed({in[726],1'b0})+$signed(in[726])+$signed(sharing147_r)+$signed(-1);
assign out[0] = (weighted_sum[0][12]==1) ? 4'd0 : (weighted_sum[0][11:8] > 6 ? 4'd6 : weighted_sum[0][11:8]);
assign out[1] = (weighted_sum[1][12]==1) ? 4'd0 : (weighted_sum[1][11:8] > 6 ? 4'd6 : weighted_sum[1][11:8]);
assign out[2] = (weighted_sum[2][12]==1) ? 4'd0 : (weighted_sum[2][11:8] > 6 ? 4'd6 : weighted_sum[2][11:8]);
assign out[3] = (weighted_sum[3][12]==1) ? 4'd0 : (weighted_sum[3][11:8] > 6 ? 4'd6 : weighted_sum[3][11:8]);
assign out[4] = (weighted_sum[4][12]==1) ? 4'd0 : (weighted_sum[4][11:8] > 6 ? 4'd6 : weighted_sum[4][11:8]);
assign out[5] = (weighted_sum[5][12]==1) ? 4'd0 : (weighted_sum[5][11:8] > 6 ? 4'd6 : weighted_sum[5][11:8]);
assign out[6] = (weighted_sum[6][12]==1) ? 4'd0 : (weighted_sum[6][11:8] > 6 ? 4'd6 : weighted_sum[6][11:8]);
assign out[7] = (weighted_sum[7][12]==1) ? 4'd0 : (weighted_sum[7][11:8] > 6 ? 4'd6 : weighted_sum[7][11:8]);
assign out[8] = (weighted_sum[8][12]==1) ? 4'd0 : (weighted_sum[8][11:8] > 6 ? 4'd6 : weighted_sum[8][11:8]);
assign out[9] = (weighted_sum[9][12]==1) ? 4'd0 : (weighted_sum[9][11:8] > 6 ? 4'd6 : weighted_sum[9][11:8]);
assign out[10] = (weighted_sum[10][12]==1) ? 4'd0 : (weighted_sum[10][11:8] > 6 ? 4'd6 : weighted_sum[10][11:8]);
assign out[11] = (weighted_sum[11][12]==1) ? 4'd0 : (weighted_sum[11][11:8] > 6 ? 4'd6 : weighted_sum[11][11:8]);
assign out[12] = (weighted_sum[12][12]==1) ? 4'd0 : (weighted_sum[12][11:8] > 6 ? 4'd6 : weighted_sum[12][11:8]);
assign out[13] = (weighted_sum[13][12]==1) ? 4'd0 : (weighted_sum[13][11:8] > 6 ? 4'd6 : weighted_sum[13][11:8]);
assign out[14] = (weighted_sum[14][12]==1) ? 4'd0 : (weighted_sum[14][11:8] > 6 ? 4'd6 : weighted_sum[14][11:8]);
assign out[15] = (weighted_sum[15][12]==1) ? 4'd0 : (weighted_sum[15][11:8] > 6 ? 4'd6 : weighted_sum[15][11:8]);
assign out[16] = (weighted_sum[16][12]==1) ? 4'd0 : (weighted_sum[16][11:8] > 6 ? 4'd6 : weighted_sum[16][11:8]);
assign out[17] = (weighted_sum[17][12]==1) ? 4'd0 : (weighted_sum[17][11:8] > 6 ? 4'd6 : weighted_sum[17][11:8]);
assign out[18] = (weighted_sum[18][12]==1) ? 4'd0 : (weighted_sum[18][11:8] > 6 ? 4'd6 : weighted_sum[18][11:8]);
assign out[19] = (weighted_sum[19][12]==1) ? 4'd0 : (weighted_sum[19][11:8] > 6 ? 4'd6 : weighted_sum[19][11:8]);
assign out[20] = (weighted_sum[20][12]==1) ? 4'd0 : (weighted_sum[20][11:8] > 6 ? 4'd6 : weighted_sum[20][11:8]);
assign out[21] = (weighted_sum[21][12]==1) ? 4'd0 : (weighted_sum[21][11:8] > 6 ? 4'd6 : weighted_sum[21][11:8]);
assign out[22] = (weighted_sum[22][12]==1) ? 4'd0 : (weighted_sum[22][11:8] > 6 ? 4'd6 : weighted_sum[22][11:8]);
assign out[23] = (weighted_sum[23][12]==1) ? 4'd0 : (weighted_sum[23][11:8] > 6 ? 4'd6 : weighted_sum[23][11:8]);
assign out[24] = (weighted_sum[24][12]==1) ? 4'd0 : (weighted_sum[24][11:8] > 6 ? 4'd6 : weighted_sum[24][11:8]);
assign out[25] = (weighted_sum[25][12]==1) ? 4'd0 : (weighted_sum[25][11:8] > 6 ? 4'd6 : weighted_sum[25][11:8]);
assign out[26] = (weighted_sum[26][12]==1) ? 4'd0 : (weighted_sum[26][11:8] > 6 ? 4'd6 : weighted_sum[26][11:8]);
assign out[27] = (weighted_sum[27][12]==1) ? 4'd0 : (weighted_sum[27][11:8] > 6 ? 4'd6 : weighted_sum[27][11:8]);
assign out[28] = (weighted_sum[28][12]==1) ? 4'd0 : (weighted_sum[28][11:8] > 6 ? 4'd6 : weighted_sum[28][11:8]);
assign out[29] = (weighted_sum[29][12]==1) ? 4'd0 : (weighted_sum[29][11:8] > 6 ? 4'd6 : weighted_sum[29][11:8]);
assign out[30] = (weighted_sum[30][12]==1) ? 4'd0 : (weighted_sum[30][11:8] > 6 ? 4'd6 : weighted_sum[30][11:8]);
assign out[31] = (weighted_sum[31][12]==1) ? 4'd0 : (weighted_sum[31][11:8] > 6 ? 4'd6 : weighted_sum[31][11:8]);
assign out[32] = (weighted_sum[32][12]==1) ? 4'd0 : (weighted_sum[32][11:8] > 6 ? 4'd6 : weighted_sum[32][11:8]);
assign out[33] = (weighted_sum[33][12]==1) ? 4'd0 : (weighted_sum[33][11:8] > 6 ? 4'd6 : weighted_sum[33][11:8]);
assign out[34] = (weighted_sum[34][12]==1) ? 4'd0 : (weighted_sum[34][11:8] > 6 ? 4'd6 : weighted_sum[34][11:8]);
assign out[35] = (weighted_sum[35][12]==1) ? 4'd0 : (weighted_sum[35][11:8] > 6 ? 4'd6 : weighted_sum[35][11:8]);
assign out[36] = (weighted_sum[36][12]==1) ? 4'd0 : (weighted_sum[36][11:8] > 6 ? 4'd6 : weighted_sum[36][11:8]);
assign out[37] = (weighted_sum[37][12]==1) ? 4'd0 : (weighted_sum[37][11:8] > 6 ? 4'd6 : weighted_sum[37][11:8]);
assign out[38] = (weighted_sum[38][12]==1) ? 4'd0 : (weighted_sum[38][11:8] > 6 ? 4'd6 : weighted_sum[38][11:8]);
assign out[39] = (weighted_sum[39][12]==1) ? 4'd0 : (weighted_sum[39][11:8] > 6 ? 4'd6 : weighted_sum[39][11:8]);
assign out[40] = (weighted_sum[40][12]==1) ? 4'd0 : (weighted_sum[40][11:8] > 6 ? 4'd6 : weighted_sum[40][11:8]);
assign out[41] = (weighted_sum[41][12]==1) ? 4'd0 : (weighted_sum[41][11:8] > 6 ? 4'd6 : weighted_sum[41][11:8]);
assign out[42] = (weighted_sum[42][12]==1) ? 4'd0 : (weighted_sum[42][11:8] > 6 ? 4'd6 : weighted_sum[42][11:8]);
assign out[43] = (weighted_sum[43][12]==1) ? 4'd0 : (weighted_sum[43][11:8] > 6 ? 4'd6 : weighted_sum[43][11:8]);
assign out[44] = (weighted_sum[44][12]==1) ? 4'd0 : (weighted_sum[44][11:8] > 6 ? 4'd6 : weighted_sum[44][11:8]);
assign out[45] = (weighted_sum[45][12]==1) ? 4'd0 : (weighted_sum[45][11:8] > 6 ? 4'd6 : weighted_sum[45][11:8]);
assign out[46] = (weighted_sum[46][12]==1) ? 4'd0 : (weighted_sum[46][11:8] > 6 ? 4'd6 : weighted_sum[46][11:8]);
assign out[47] = (weighted_sum[47][12]==1) ? 4'd0 : (weighted_sum[47][11:8] > 6 ? 4'd6 : weighted_sum[47][11:8]);
assign out[48] = (weighted_sum[48][12]==1) ? 4'd0 : (weighted_sum[48][11:8] > 6 ? 4'd6 : weighted_sum[48][11:8]);
assign out[49] = (weighted_sum[49][12]==1) ? 4'd0 : (weighted_sum[49][11:8] > 6 ? 4'd6 : weighted_sum[49][11:8]);
assign out[50] = (weighted_sum[50][12]==1) ? 4'd0 : (weighted_sum[50][11:8] > 6 ? 4'd6 : weighted_sum[50][11:8]);
assign out[51] = (weighted_sum[51][12]==1) ? 4'd0 : (weighted_sum[51][11:8] > 6 ? 4'd6 : weighted_sum[51][11:8]);
assign out[52] = (weighted_sum[52][12]==1) ? 4'd0 : (weighted_sum[52][11:8] > 6 ? 4'd6 : weighted_sum[52][11:8]);
assign out[53] = (weighted_sum[53][12]==1) ? 4'd0 : (weighted_sum[53][11:8] > 6 ? 4'd6 : weighted_sum[53][11:8]);
assign out[54] = (weighted_sum[54][12]==1) ? 4'd0 : (weighted_sum[54][11:8] > 6 ? 4'd6 : weighted_sum[54][11:8]);
assign out[55] = (weighted_sum[55][12]==1) ? 4'd0 : (weighted_sum[55][11:8] > 6 ? 4'd6 : weighted_sum[55][11:8]);
assign out[56] = (weighted_sum[56][12]==1) ? 4'd0 : (weighted_sum[56][11:8] > 6 ? 4'd6 : weighted_sum[56][11:8]);
assign out[57] = (weighted_sum[57][12]==1) ? 4'd0 : (weighted_sum[57][11:8] > 6 ? 4'd6 : weighted_sum[57][11:8]);
assign out[58] = (weighted_sum[58][12]==1) ? 4'd0 : (weighted_sum[58][11:8] > 6 ? 4'd6 : weighted_sum[58][11:8]);
assign out[59] = (weighted_sum[59][12]==1) ? 4'd0 : (weighted_sum[59][11:8] > 6 ? 4'd6 : weighted_sum[59][11:8]);
assign out[60] = (weighted_sum[60][12]==1) ? 4'd0 : (weighted_sum[60][11:8] > 6 ? 4'd6 : weighted_sum[60][11:8]);
assign out[61] = (weighted_sum[61][12]==1) ? 4'd0 : (weighted_sum[61][11:8] > 6 ? 4'd6 : weighted_sum[61][11:8]);
assign out[62] = (weighted_sum[62][12]==1) ? 4'd0 : (weighted_sum[62][11:8] > 6 ? 4'd6 : weighted_sum[62][11:8]);
assign out[63] = (weighted_sum[63][12]==1) ? 4'd0 : (weighted_sum[63][11:8] > 6 ? 4'd6 : weighted_sum[63][11:8]);
assign out[64] = (weighted_sum[64][12]==1) ? 4'd0 : (weighted_sum[64][11:8] > 6 ? 4'd6 : weighted_sum[64][11:8]);
assign out[65] = (weighted_sum[65][12]==1) ? 4'd0 : (weighted_sum[65][11:8] > 6 ? 4'd6 : weighted_sum[65][11:8]);
assign out[66] = (weighted_sum[66][12]==1) ? 4'd0 : (weighted_sum[66][11:8] > 6 ? 4'd6 : weighted_sum[66][11:8]);
assign out[67] = (weighted_sum[67][12]==1) ? 4'd0 : (weighted_sum[67][11:8] > 6 ? 4'd6 : weighted_sum[67][11:8]);
assign out[68] = (weighted_sum[68][12]==1) ? 4'd0 : (weighted_sum[68][11:8] > 6 ? 4'd6 : weighted_sum[68][11:8]);
assign out[69] = (weighted_sum[69][12]==1) ? 4'd0 : (weighted_sum[69][11:8] > 6 ? 4'd6 : weighted_sum[69][11:8]);
assign out[70] = (weighted_sum[70][12]==1) ? 4'd0 : (weighted_sum[70][11:8] > 6 ? 4'd6 : weighted_sum[70][11:8]);
assign out[71] = (weighted_sum[71][12]==1) ? 4'd0 : (weighted_sum[71][11:8] > 6 ? 4'd6 : weighted_sum[71][11:8]);
assign out[72] = (weighted_sum[72][12]==1) ? 4'd0 : (weighted_sum[72][11:8] > 6 ? 4'd6 : weighted_sum[72][11:8]);
assign out[73] = (weighted_sum[73][12]==1) ? 4'd0 : (weighted_sum[73][11:8] > 6 ? 4'd6 : weighted_sum[73][11:8]);
assign out[74] = (weighted_sum[74][12]==1) ? 4'd0 : (weighted_sum[74][11:8] > 6 ? 4'd6 : weighted_sum[74][11:8]);
assign out[75] = (weighted_sum[75][12]==1) ? 4'd0 : (weighted_sum[75][11:8] > 6 ? 4'd6 : weighted_sum[75][11:8]);
assign out[76] = (weighted_sum[76][12]==1) ? 4'd0 : (weighted_sum[76][11:8] > 6 ? 4'd6 : weighted_sum[76][11:8]);
assign out[77] = (weighted_sum[77][12]==1) ? 4'd0 : (weighted_sum[77][11:8] > 6 ? 4'd6 : weighted_sum[77][11:8]);
assign out[78] = (weighted_sum[78][12]==1) ? 4'd0 : (weighted_sum[78][11:8] > 6 ? 4'd6 : weighted_sum[78][11:8]);
assign out[79] = (weighted_sum[79][12]==1) ? 4'd0 : (weighted_sum[79][11:8] > 6 ? 4'd6 : weighted_sum[79][11:8]);
assign out[80] = (weighted_sum[80][12]==1) ? 4'd0 : (weighted_sum[80][11:8] > 6 ? 4'd6 : weighted_sum[80][11:8]);
assign out[81] = (weighted_sum[81][12]==1) ? 4'd0 : (weighted_sum[81][11:8] > 6 ? 4'd6 : weighted_sum[81][11:8]);
assign out[82] = (weighted_sum[82][12]==1) ? 4'd0 : (weighted_sum[82][11:8] > 6 ? 4'd6 : weighted_sum[82][11:8]);
assign out[83] = (weighted_sum[83][12]==1) ? 4'd0 : (weighted_sum[83][11:8] > 6 ? 4'd6 : weighted_sum[83][11:8]);
assign out[84] = (weighted_sum[84][12]==1) ? 4'd0 : (weighted_sum[84][11:8] > 6 ? 4'd6 : weighted_sum[84][11:8]);
assign out[85] = (weighted_sum[85][12]==1) ? 4'd0 : (weighted_sum[85][11:8] > 6 ? 4'd6 : weighted_sum[85][11:8]);
assign out[86] = (weighted_sum[86][12]==1) ? 4'd0 : (weighted_sum[86][11:8] > 6 ? 4'd6 : weighted_sum[86][11:8]);
assign out[87] = (weighted_sum[87][12]==1) ? 4'd0 : (weighted_sum[87][11:8] > 6 ? 4'd6 : weighted_sum[87][11:8]);
assign out[88] = (weighted_sum[88][12]==1) ? 4'd0 : (weighted_sum[88][11:8] > 6 ? 4'd6 : weighted_sum[88][11:8]);
assign out[89] = (weighted_sum[89][12]==1) ? 4'd0 : (weighted_sum[89][11:8] > 6 ? 4'd6 : weighted_sum[89][11:8]);
assign out[90] = (weighted_sum[90][12]==1) ? 4'd0 : (weighted_sum[90][11:8] > 6 ? 4'd6 : weighted_sum[90][11:8]);
assign out[91] = (weighted_sum[91][12]==1) ? 4'd0 : (weighted_sum[91][11:8] > 6 ? 4'd6 : weighted_sum[91][11:8]);
assign out[92] = (weighted_sum[92][12]==1) ? 4'd0 : (weighted_sum[92][11:8] > 6 ? 4'd6 : weighted_sum[92][11:8]);
assign out[93] = (weighted_sum[93][12]==1) ? 4'd0 : (weighted_sum[93][11:8] > 6 ? 4'd6 : weighted_sum[93][11:8]);
assign out[94] = (weighted_sum[94][12]==1) ? 4'd0 : (weighted_sum[94][11:8] > 6 ? 4'd6 : weighted_sum[94][11:8]);
assign out[95] = (weighted_sum[95][12]==1) ? 4'd0 : (weighted_sum[95][11:8] > 6 ? 4'd6 : weighted_sum[95][11:8]);
assign out[96] = (weighted_sum[96][12]==1) ? 4'd0 : (weighted_sum[96][11:8] > 6 ? 4'd6 : weighted_sum[96][11:8]);
assign out[97] = (weighted_sum[97][12]==1) ? 4'd0 : (weighted_sum[97][11:8] > 6 ? 4'd6 : weighted_sum[97][11:8]);
assign out[98] = (weighted_sum[98][12]==1) ? 4'd0 : (weighted_sum[98][11:8] > 6 ? 4'd6 : weighted_sum[98][11:8]);
assign out[99] = (weighted_sum[99][12]==1) ? 4'd0 : (weighted_sum[99][11:8] > 6 ? 4'd6 : weighted_sum[99][11:8]);
assign out[100] = (weighted_sum[100][12]==1) ? 4'd0 : (weighted_sum[100][11:8] > 6 ? 4'd6 : weighted_sum[100][11:8]);
assign out[101] = (weighted_sum[101][12]==1) ? 4'd0 : (weighted_sum[101][11:8] > 6 ? 4'd6 : weighted_sum[101][11:8]);
assign out[102] = (weighted_sum[102][12]==1) ? 4'd0 : (weighted_sum[102][11:8] > 6 ? 4'd6 : weighted_sum[102][11:8]);
assign out[103] = (weighted_sum[103][12]==1) ? 4'd0 : (weighted_sum[103][11:8] > 6 ? 4'd6 : weighted_sum[103][11:8]);
assign out[104] = (weighted_sum[104][12]==1) ? 4'd0 : (weighted_sum[104][11:8] > 6 ? 4'd6 : weighted_sum[104][11:8]);
assign out[105] = (weighted_sum[105][12]==1) ? 4'd0 : (weighted_sum[105][11:8] > 6 ? 4'd6 : weighted_sum[105][11:8]);
assign out[106] = (weighted_sum[106][12]==1) ? 4'd0 : (weighted_sum[106][11:8] > 6 ? 4'd6 : weighted_sum[106][11:8]);
assign out[107] = (weighted_sum[107][12]==1) ? 4'd0 : (weighted_sum[107][11:8] > 6 ? 4'd6 : weighted_sum[107][11:8]);
assign out[108] = (weighted_sum[108][12]==1) ? 4'd0 : (weighted_sum[108][11:8] > 6 ? 4'd6 : weighted_sum[108][11:8]);
assign out[109] = (weighted_sum[109][12]==1) ? 4'd0 : (weighted_sum[109][11:8] > 6 ? 4'd6 : weighted_sum[109][11:8]);
assign out[110] = (weighted_sum[110][12]==1) ? 4'd0 : (weighted_sum[110][11:8] > 6 ? 4'd6 : weighted_sum[110][11:8]);
assign out[111] = (weighted_sum[111][12]==1) ? 4'd0 : (weighted_sum[111][11:8] > 6 ? 4'd6 : weighted_sum[111][11:8]);
assign out[112] = (weighted_sum[112][12]==1) ? 4'd0 : (weighted_sum[112][11:8] > 6 ? 4'd6 : weighted_sum[112][11:8]);
assign out[113] = (weighted_sum[113][12]==1) ? 4'd0 : (weighted_sum[113][11:8] > 6 ? 4'd6 : weighted_sum[113][11:8]);
assign out[114] = (weighted_sum[114][12]==1) ? 4'd0 : (weighted_sum[114][11:8] > 6 ? 4'd6 : weighted_sum[114][11:8]);
assign out[115] = (weighted_sum[115][12]==1) ? 4'd0 : (weighted_sum[115][11:8] > 6 ? 4'd6 : weighted_sum[115][11:8]);
assign out[116] = (weighted_sum[116][12]==1) ? 4'd0 : (weighted_sum[116][11:8] > 6 ? 4'd6 : weighted_sum[116][11:8]);
assign out[117] = (weighted_sum[117][12]==1) ? 4'd0 : (weighted_sum[117][11:8] > 6 ? 4'd6 : weighted_sum[117][11:8]);
assign out[118] = (weighted_sum[118][12]==1) ? 4'd0 : (weighted_sum[118][11:8] > 6 ? 4'd6 : weighted_sum[118][11:8]);
assign out[119] = (weighted_sum[119][12]==1) ? 4'd0 : (weighted_sum[119][11:8] > 6 ? 4'd6 : weighted_sum[119][11:8]);
assign out[120] = (weighted_sum[120][12]==1) ? 4'd0 : (weighted_sum[120][11:8] > 6 ? 4'd6 : weighted_sum[120][11:8]);
assign out[121] = (weighted_sum[121][12]==1) ? 4'd0 : (weighted_sum[121][11:8] > 6 ? 4'd6 : weighted_sum[121][11:8]);
assign out[122] = (weighted_sum[122][12]==1) ? 4'd0 : (weighted_sum[122][11:8] > 6 ? 4'd6 : weighted_sum[122][11:8]);
assign out[123] = (weighted_sum[123][12]==1) ? 4'd0 : (weighted_sum[123][11:8] > 6 ? 4'd6 : weighted_sum[123][11:8]);
assign out[124] = (weighted_sum[124][12]==1) ? 4'd0 : (weighted_sum[124][11:8] > 6 ? 4'd6 : weighted_sum[124][11:8]);
assign out[125] = (weighted_sum[125][12]==1) ? 4'd0 : (weighted_sum[125][11:8] > 6 ? 4'd6 : weighted_sum[125][11:8]);
assign out[126] = (weighted_sum[126][12]==1) ? 4'd0 : (weighted_sum[126][11:8] > 6 ? 4'd6 : weighted_sum[126][11:8]);
assign out[127] = (weighted_sum[127][12]==1) ? 4'd0 : (weighted_sum[127][11:8] > 6 ? 4'd6 : weighted_sum[127][11:8]);
assign out[128] = (weighted_sum[128][12]==1) ? 4'd0 : (weighted_sum[128][11:8] > 6 ? 4'd6 : weighted_sum[128][11:8]);
assign out[129] = (weighted_sum[129][12]==1) ? 4'd0 : (weighted_sum[129][11:8] > 6 ? 4'd6 : weighted_sum[129][11:8]);
assign out[130] = (weighted_sum[130][12]==1) ? 4'd0 : (weighted_sum[130][11:8] > 6 ? 4'd6 : weighted_sum[130][11:8]);
assign out[131] = (weighted_sum[131][12]==1) ? 4'd0 : (weighted_sum[131][11:8] > 6 ? 4'd6 : weighted_sum[131][11:8]);
assign out[132] = (weighted_sum[132][12]==1) ? 4'd0 : (weighted_sum[132][11:8] > 6 ? 4'd6 : weighted_sum[132][11:8]);
assign out[133] = (weighted_sum[133][12]==1) ? 4'd0 : (weighted_sum[133][11:8] > 6 ? 4'd6 : weighted_sum[133][11:8]);
assign out[134] = (weighted_sum[134][12]==1) ? 4'd0 : (weighted_sum[134][11:8] > 6 ? 4'd6 : weighted_sum[134][11:8]);
assign out[135] = (weighted_sum[135][12]==1) ? 4'd0 : (weighted_sum[135][11:8] > 6 ? 4'd6 : weighted_sum[135][11:8]);
assign out[136] = (weighted_sum[136][12]==1) ? 4'd0 : (weighted_sum[136][11:8] > 6 ? 4'd6 : weighted_sum[136][11:8]);
assign out[137] = (weighted_sum[137][12]==1) ? 4'd0 : (weighted_sum[137][11:8] > 6 ? 4'd6 : weighted_sum[137][11:8]);
assign out[138] = (weighted_sum[138][12]==1) ? 4'd0 : (weighted_sum[138][11:8] > 6 ? 4'd6 : weighted_sum[138][11:8]);
assign out[139] = (weighted_sum[139][12]==1) ? 4'd0 : (weighted_sum[139][11:8] > 6 ? 4'd6 : weighted_sum[139][11:8]);
assign out[140] = (weighted_sum[140][12]==1) ? 4'd0 : (weighted_sum[140][11:8] > 6 ? 4'd6 : weighted_sum[140][11:8]);
assign out[141] = (weighted_sum[141][12]==1) ? 4'd0 : (weighted_sum[141][11:8] > 6 ? 4'd6 : weighted_sum[141][11:8]);
assign out[142] = (weighted_sum[142][12]==1) ? 4'd0 : (weighted_sum[142][11:8] > 6 ? 4'd6 : weighted_sum[142][11:8]);
assign out[143] = (weighted_sum[143][12]==1) ? 4'd0 : (weighted_sum[143][11:8] > 6 ? 4'd6 : weighted_sum[143][11:8]);
assign out[144] = (weighted_sum[144][12]==1) ? 4'd0 : (weighted_sum[144][11:8] > 6 ? 4'd6 : weighted_sum[144][11:8]);
assign out[145] = (weighted_sum[145][12]==1) ? 4'd0 : (weighted_sum[145][11:8] > 6 ? 4'd6 : weighted_sum[145][11:8]);
assign out[146] = (weighted_sum[146][12]==1) ? 4'd0 : (weighted_sum[146][11:8] > 6 ? 4'd6 : weighted_sum[146][11:8]);
assign out[147] = (weighted_sum[147][12]==1) ? 4'd0 : (weighted_sum[147][11:8] > 6 ? 4'd6 : weighted_sum[147][11:8]);
assign out[148] = (weighted_sum[148][12]==1) ? 4'd0 : (weighted_sum[148][11:8] > 6 ? 4'd6 : weighted_sum[148][11:8]);
assign out[149] = (weighted_sum[149][12]==1) ? 4'd0 : (weighted_sum[149][11:8] > 6 ? 4'd6 : weighted_sum[149][11:8]);
assign out[150] = (weighted_sum[150][12]==1) ? 4'd0 : (weighted_sum[150][11:8] > 6 ? 4'd6 : weighted_sum[150][11:8]);
assign out[151] = (weighted_sum[151][12]==1) ? 4'd0 : (weighted_sum[151][11:8] > 6 ? 4'd6 : weighted_sum[151][11:8]);
assign out[152] = (weighted_sum[152][12]==1) ? 4'd0 : (weighted_sum[152][11:8] > 6 ? 4'd6 : weighted_sum[152][11:8]);
assign out[153] = (weighted_sum[153][12]==1) ? 4'd0 : (weighted_sum[153][11:8] > 6 ? 4'd6 : weighted_sum[153][11:8]);
assign out[154] = (weighted_sum[154][12]==1) ? 4'd0 : (weighted_sum[154][11:8] > 6 ? 4'd6 : weighted_sum[154][11:8]);
assign out[155] = (weighted_sum[155][12]==1) ? 4'd0 : (weighted_sum[155][11:8] > 6 ? 4'd6 : weighted_sum[155][11:8]);
assign out[156] = (weighted_sum[156][12]==1) ? 4'd0 : (weighted_sum[156][11:8] > 6 ? 4'd6 : weighted_sum[156][11:8]);
assign out[157] = (weighted_sum[157][12]==1) ? 4'd0 : (weighted_sum[157][11:8] > 6 ? 4'd6 : weighted_sum[157][11:8]);
assign out[158] = (weighted_sum[158][12]==1) ? 4'd0 : (weighted_sum[158][11:8] > 6 ? 4'd6 : weighted_sum[158][11:8]);
assign out[159] = (weighted_sum[159][12]==1) ? 4'd0 : (weighted_sum[159][11:8] > 6 ? 4'd6 : weighted_sum[159][11:8]);
assign out[160] = (weighted_sum[160][12]==1) ? 4'd0 : (weighted_sum[160][11:8] > 6 ? 4'd6 : weighted_sum[160][11:8]);
assign out[161] = (weighted_sum[161][12]==1) ? 4'd0 : (weighted_sum[161][11:8] > 6 ? 4'd6 : weighted_sum[161][11:8]);
assign out[162] = (weighted_sum[162][12]==1) ? 4'd0 : (weighted_sum[162][11:8] > 6 ? 4'd6 : weighted_sum[162][11:8]);
assign out[163] = (weighted_sum[163][12]==1) ? 4'd0 : (weighted_sum[163][11:8] > 6 ? 4'd6 : weighted_sum[163][11:8]);
assign out[164] = (weighted_sum[164][12]==1) ? 4'd0 : (weighted_sum[164][11:8] > 6 ? 4'd6 : weighted_sum[164][11:8]);
assign out[165] = (weighted_sum[165][12]==1) ? 4'd0 : (weighted_sum[165][11:8] > 6 ? 4'd6 : weighted_sum[165][11:8]);
assign out[166] = (weighted_sum[166][12]==1) ? 4'd0 : (weighted_sum[166][11:8] > 6 ? 4'd6 : weighted_sum[166][11:8]);
assign out[167] = (weighted_sum[167][12]==1) ? 4'd0 : (weighted_sum[167][11:8] > 6 ? 4'd6 : weighted_sum[167][11:8]);
assign out[168] = (weighted_sum[168][12]==1) ? 4'd0 : (weighted_sum[168][11:8] > 6 ? 4'd6 : weighted_sum[168][11:8]);
assign out[169] = (weighted_sum[169][12]==1) ? 4'd0 : (weighted_sum[169][11:8] > 6 ? 4'd6 : weighted_sum[169][11:8]);
assign out[170] = (weighted_sum[170][12]==1) ? 4'd0 : (weighted_sum[170][11:8] > 6 ? 4'd6 : weighted_sum[170][11:8]);
assign out[171] = (weighted_sum[171][12]==1) ? 4'd0 : (weighted_sum[171][11:8] > 6 ? 4'd6 : weighted_sum[171][11:8]);
assign out[172] = (weighted_sum[172][12]==1) ? 4'd0 : (weighted_sum[172][11:8] > 6 ? 4'd6 : weighted_sum[172][11:8]);
assign out[173] = (weighted_sum[173][12]==1) ? 4'd0 : (weighted_sum[173][11:8] > 6 ? 4'd6 : weighted_sum[173][11:8]);
assign out[174] = (weighted_sum[174][12]==1) ? 4'd0 : (weighted_sum[174][11:8] > 6 ? 4'd6 : weighted_sum[174][11:8]);
assign out[175] = (weighted_sum[175][12]==1) ? 4'd0 : (weighted_sum[175][11:8] > 6 ? 4'd6 : weighted_sum[175][11:8]);
assign out[176] = (weighted_sum[176][12]==1) ? 4'd0 : (weighted_sum[176][11:8] > 6 ? 4'd6 : weighted_sum[176][11:8]);
assign out[177] = (weighted_sum[177][12]==1) ? 4'd0 : (weighted_sum[177][11:8] > 6 ? 4'd6 : weighted_sum[177][11:8]);
assign out[178] = (weighted_sum[178][12]==1) ? 4'd0 : (weighted_sum[178][11:8] > 6 ? 4'd6 : weighted_sum[178][11:8]);
assign out[179] = (weighted_sum[179][12]==1) ? 4'd0 : (weighted_sum[179][11:8] > 6 ? 4'd6 : weighted_sum[179][11:8]);
assign out[180] = (weighted_sum[180][12]==1) ? 4'd0 : (weighted_sum[180][11:8] > 6 ? 4'd6 : weighted_sum[180][11:8]);
assign out[181] = (weighted_sum[181][12]==1) ? 4'd0 : (weighted_sum[181][11:8] > 6 ? 4'd6 : weighted_sum[181][11:8]);
assign out[182] = (weighted_sum[182][12]==1) ? 4'd0 : (weighted_sum[182][11:8] > 6 ? 4'd6 : weighted_sum[182][11:8]);
assign out[183] = (weighted_sum[183][12]==1) ? 4'd0 : (weighted_sum[183][11:8] > 6 ? 4'd6 : weighted_sum[183][11:8]);
assign out[184] = (weighted_sum[184][12]==1) ? 4'd0 : (weighted_sum[184][11:8] > 6 ? 4'd6 : weighted_sum[184][11:8]);
assign out[185] = (weighted_sum[185][12]==1) ? 4'd0 : (weighted_sum[185][11:8] > 6 ? 4'd6 : weighted_sum[185][11:8]);
assign out[186] = (weighted_sum[186][12]==1) ? 4'd0 : (weighted_sum[186][11:8] > 6 ? 4'd6 : weighted_sum[186][11:8]);
assign out[187] = (weighted_sum[187][12]==1) ? 4'd0 : (weighted_sum[187][11:8] > 6 ? 4'd6 : weighted_sum[187][11:8]);
assign out[188] = (weighted_sum[188][12]==1) ? 4'd0 : (weighted_sum[188][11:8] > 6 ? 4'd6 : weighted_sum[188][11:8]);
assign out[189] = (weighted_sum[189][12]==1) ? 4'd0 : (weighted_sum[189][11:8] > 6 ? 4'd6 : weighted_sum[189][11:8]);
assign out[190] = (weighted_sum[190][12]==1) ? 4'd0 : (weighted_sum[190][11:8] > 6 ? 4'd6 : weighted_sum[190][11:8]);
assign out[191] = (weighted_sum[191][12]==1) ? 4'd0 : (weighted_sum[191][11:8] > 6 ? 4'd6 : weighted_sum[191][11:8]);
assign out[192] = (weighted_sum[192][12]==1) ? 4'd0 : (weighted_sum[192][11:8] > 6 ? 4'd6 : weighted_sum[192][11:8]);
assign out[193] = (weighted_sum[193][12]==1) ? 4'd0 : (weighted_sum[193][11:8] > 6 ? 4'd6 : weighted_sum[193][11:8]);
assign out[194] = (weighted_sum[194][12]==1) ? 4'd0 : (weighted_sum[194][11:8] > 6 ? 4'd6 : weighted_sum[194][11:8]);
assign out[195] = (weighted_sum[195][12]==1) ? 4'd0 : (weighted_sum[195][11:8] > 6 ? 4'd6 : weighted_sum[195][11:8]);
assign out[196] = (weighted_sum[196][12]==1) ? 4'd0 : (weighted_sum[196][11:8] > 6 ? 4'd6 : weighted_sum[196][11:8]);
assign out[197] = (weighted_sum[197][12]==1) ? 4'd0 : (weighted_sum[197][11:8] > 6 ? 4'd6 : weighted_sum[197][11:8]);
assign out[198] = (weighted_sum[198][12]==1) ? 4'd0 : (weighted_sum[198][11:8] > 6 ? 4'd6 : weighted_sum[198][11:8]);
assign out[199] = (weighted_sum[199][12]==1) ? 4'd0 : (weighted_sum[199][11:8] > 6 ? 4'd6 : weighted_sum[199][11:8]);
assign out[200] = (weighted_sum[200][12]==1) ? 4'd0 : (weighted_sum[200][11:8] > 6 ? 4'd6 : weighted_sum[200][11:8]);
assign out[201] = (weighted_sum[201][12]==1) ? 4'd0 : (weighted_sum[201][11:8] > 6 ? 4'd6 : weighted_sum[201][11:8]);
assign out[202] = (weighted_sum[202][12]==1) ? 4'd0 : (weighted_sum[202][11:8] > 6 ? 4'd6 : weighted_sum[202][11:8]);
assign out[203] = (weighted_sum[203][12]==1) ? 4'd0 : (weighted_sum[203][11:8] > 6 ? 4'd6 : weighted_sum[203][11:8]);
assign out[204] = (weighted_sum[204][12]==1) ? 4'd0 : (weighted_sum[204][11:8] > 6 ? 4'd6 : weighted_sum[204][11:8]);
assign out[205] = (weighted_sum[205][12]==1) ? 4'd0 : (weighted_sum[205][11:8] > 6 ? 4'd6 : weighted_sum[205][11:8]);
assign out[206] = (weighted_sum[206][12]==1) ? 4'd0 : (weighted_sum[206][11:8] > 6 ? 4'd6 : weighted_sum[206][11:8]);
assign out[207] = (weighted_sum[207][12]==1) ? 4'd0 : (weighted_sum[207][11:8] > 6 ? 4'd6 : weighted_sum[207][11:8]);
assign out[208] = (weighted_sum[208][12]==1) ? 4'd0 : (weighted_sum[208][11:8] > 6 ? 4'd6 : weighted_sum[208][11:8]);
assign out[209] = (weighted_sum[209][12]==1) ? 4'd0 : (weighted_sum[209][11:8] > 6 ? 4'd6 : weighted_sum[209][11:8]);
assign out[210] = (weighted_sum[210][12]==1) ? 4'd0 : (weighted_sum[210][11:8] > 6 ? 4'd6 : weighted_sum[210][11:8]);
assign out[211] = (weighted_sum[211][12]==1) ? 4'd0 : (weighted_sum[211][11:8] > 6 ? 4'd6 : weighted_sum[211][11:8]);
assign out[212] = (weighted_sum[212][12]==1) ? 4'd0 : (weighted_sum[212][11:8] > 6 ? 4'd6 : weighted_sum[212][11:8]);
assign out[213] = (weighted_sum[213][12]==1) ? 4'd0 : (weighted_sum[213][11:8] > 6 ? 4'd6 : weighted_sum[213][11:8]);
assign out[214] = (weighted_sum[214][12]==1) ? 4'd0 : (weighted_sum[214][11:8] > 6 ? 4'd6 : weighted_sum[214][11:8]);
assign out[215] = (weighted_sum[215][12]==1) ? 4'd0 : (weighted_sum[215][11:8] > 6 ? 4'd6 : weighted_sum[215][11:8]);
assign out[216] = (weighted_sum[216][12]==1) ? 4'd0 : (weighted_sum[216][11:8] > 6 ? 4'd6 : weighted_sum[216][11:8]);
assign out[217] = (weighted_sum[217][12]==1) ? 4'd0 : (weighted_sum[217][11:8] > 6 ? 4'd6 : weighted_sum[217][11:8]);
assign out[218] = (weighted_sum[218][12]==1) ? 4'd0 : (weighted_sum[218][11:8] > 6 ? 4'd6 : weighted_sum[218][11:8]);
assign out[219] = (weighted_sum[219][12]==1) ? 4'd0 : (weighted_sum[219][11:8] > 6 ? 4'd6 : weighted_sum[219][11:8]);
assign out[220] = (weighted_sum[220][12]==1) ? 4'd0 : (weighted_sum[220][11:8] > 6 ? 4'd6 : weighted_sum[220][11:8]);
assign out[221] = (weighted_sum[221][12]==1) ? 4'd0 : (weighted_sum[221][11:8] > 6 ? 4'd6 : weighted_sum[221][11:8]);
assign out[222] = (weighted_sum[222][12]==1) ? 4'd0 : (weighted_sum[222][11:8] > 6 ? 4'd6 : weighted_sum[222][11:8]);
assign out[223] = (weighted_sum[223][12]==1) ? 4'd0 : (weighted_sum[223][11:8] > 6 ? 4'd6 : weighted_sum[223][11:8]);
assign out[224] = (weighted_sum[224][12]==1) ? 4'd0 : (weighted_sum[224][11:8] > 6 ? 4'd6 : weighted_sum[224][11:8]);
assign out[225] = (weighted_sum[225][12]==1) ? 4'd0 : (weighted_sum[225][11:8] > 6 ? 4'd6 : weighted_sum[225][11:8]);
assign out[226] = (weighted_sum[226][12]==1) ? 4'd0 : (weighted_sum[226][11:8] > 6 ? 4'd6 : weighted_sum[226][11:8]);
assign out[227] = (weighted_sum[227][12]==1) ? 4'd0 : (weighted_sum[227][11:8] > 6 ? 4'd6 : weighted_sum[227][11:8]);
assign out[228] = (weighted_sum[228][12]==1) ? 4'd0 : (weighted_sum[228][11:8] > 6 ? 4'd6 : weighted_sum[228][11:8]);
assign out[229] = (weighted_sum[229][12]==1) ? 4'd0 : (weighted_sum[229][11:8] > 6 ? 4'd6 : weighted_sum[229][11:8]);
assign out[230] = (weighted_sum[230][12]==1) ? 4'd0 : (weighted_sum[230][11:8] > 6 ? 4'd6 : weighted_sum[230][11:8]);
assign out[231] = (weighted_sum[231][12]==1) ? 4'd0 : (weighted_sum[231][11:8] > 6 ? 4'd6 : weighted_sum[231][11:8]);
assign out[232] = (weighted_sum[232][12]==1) ? 4'd0 : (weighted_sum[232][11:8] > 6 ? 4'd6 : weighted_sum[232][11:8]);
assign out[233] = (weighted_sum[233][12]==1) ? 4'd0 : (weighted_sum[233][11:8] > 6 ? 4'd6 : weighted_sum[233][11:8]);
assign out[234] = (weighted_sum[234][12]==1) ? 4'd0 : (weighted_sum[234][11:8] > 6 ? 4'd6 : weighted_sum[234][11:8]);
assign out[235] = (weighted_sum[235][12]==1) ? 4'd0 : (weighted_sum[235][11:8] > 6 ? 4'd6 : weighted_sum[235][11:8]);
assign out[236] = (weighted_sum[236][12]==1) ? 4'd0 : (weighted_sum[236][11:8] > 6 ? 4'd6 : weighted_sum[236][11:8]);
assign out[237] = (weighted_sum[237][12]==1) ? 4'd0 : (weighted_sum[237][11:8] > 6 ? 4'd6 : weighted_sum[237][11:8]);
assign out[238] = (weighted_sum[238][12]==1) ? 4'd0 : (weighted_sum[238][11:8] > 6 ? 4'd6 : weighted_sum[238][11:8]);
assign out[239] = (weighted_sum[239][12]==1) ? 4'd0 : (weighted_sum[239][11:8] > 6 ? 4'd6 : weighted_sum[239][11:8]);
assign out[240] = (weighted_sum[240][12]==1) ? 4'd0 : (weighted_sum[240][11:8] > 6 ? 4'd6 : weighted_sum[240][11:8]);
assign out[241] = (weighted_sum[241][12]==1) ? 4'd0 : (weighted_sum[241][11:8] > 6 ? 4'd6 : weighted_sum[241][11:8]);
assign out[242] = (weighted_sum[242][12]==1) ? 4'd0 : (weighted_sum[242][11:8] > 6 ? 4'd6 : weighted_sum[242][11:8]);
assign out[243] = (weighted_sum[243][12]==1) ? 4'd0 : (weighted_sum[243][11:8] > 6 ? 4'd6 : weighted_sum[243][11:8]);
assign out[244] = (weighted_sum[244][12]==1) ? 4'd0 : (weighted_sum[244][11:8] > 6 ? 4'd6 : weighted_sum[244][11:8]);
assign out[245] = (weighted_sum[245][12]==1) ? 4'd0 : (weighted_sum[245][11:8] > 6 ? 4'd6 : weighted_sum[245][11:8]);
assign out[246] = (weighted_sum[246][12]==1) ? 4'd0 : (weighted_sum[246][11:8] > 6 ? 4'd6 : weighted_sum[246][11:8]);
assign out[247] = (weighted_sum[247][12]==1) ? 4'd0 : (weighted_sum[247][11:8] > 6 ? 4'd6 : weighted_sum[247][11:8]);
assign out[248] = (weighted_sum[248][12]==1) ? 4'd0 : (weighted_sum[248][11:8] > 6 ? 4'd6 : weighted_sum[248][11:8]);
assign out[249] = (weighted_sum[249][12]==1) ? 4'd0 : (weighted_sum[249][11:8] > 6 ? 4'd6 : weighted_sum[249][11:8]);
assign out[250] = (weighted_sum[250][12]==1) ? 4'd0 : (weighted_sum[250][11:8] > 6 ? 4'd6 : weighted_sum[250][11:8]);
assign out[251] = (weighted_sum[251][12]==1) ? 4'd0 : (weighted_sum[251][11:8] > 6 ? 4'd6 : weighted_sum[251][11:8]);
assign out[252] = (weighted_sum[252][12]==1) ? 4'd0 : (weighted_sum[252][11:8] > 6 ? 4'd6 : weighted_sum[252][11:8]);
assign out[253] = (weighted_sum[253][12]==1) ? 4'd0 : (weighted_sum[253][11:8] > 6 ? 4'd6 : weighted_sum[253][11:8]);
assign out[254] = (weighted_sum[254][12]==1) ? 4'd0 : (weighted_sum[254][11:8] > 6 ? 4'd6 : weighted_sum[254][11:8]);
assign out[255] = (weighted_sum[255][12]==1) ? 4'd0 : (weighted_sum[255][11:8] > 6 ? 4'd6 : weighted_sum[255][11:8]);
assign out[256] = (weighted_sum[256][12]==1) ? 4'd0 : (weighted_sum[256][11:8] > 6 ? 4'd6 : weighted_sum[256][11:8]);
assign out[257] = (weighted_sum[257][12]==1) ? 4'd0 : (weighted_sum[257][11:8] > 6 ? 4'd6 : weighted_sum[257][11:8]);
assign out[258] = (weighted_sum[258][12]==1) ? 4'd0 : (weighted_sum[258][11:8] > 6 ? 4'd6 : weighted_sum[258][11:8]);
assign out[259] = (weighted_sum[259][12]==1) ? 4'd0 : (weighted_sum[259][11:8] > 6 ? 4'd6 : weighted_sum[259][11:8]);
assign out[260] = (weighted_sum[260][12]==1) ? 4'd0 : (weighted_sum[260][11:8] > 6 ? 4'd6 : weighted_sum[260][11:8]);
assign out[261] = (weighted_sum[261][12]==1) ? 4'd0 : (weighted_sum[261][11:8] > 6 ? 4'd6 : weighted_sum[261][11:8]);
assign out[262] = (weighted_sum[262][12]==1) ? 4'd0 : (weighted_sum[262][11:8] > 6 ? 4'd6 : weighted_sum[262][11:8]);
assign out[263] = (weighted_sum[263][12]==1) ? 4'd0 : (weighted_sum[263][11:8] > 6 ? 4'd6 : weighted_sum[263][11:8]);
assign out[264] = (weighted_sum[264][12]==1) ? 4'd0 : (weighted_sum[264][11:8] > 6 ? 4'd6 : weighted_sum[264][11:8]);
assign out[265] = (weighted_sum[265][12]==1) ? 4'd0 : (weighted_sum[265][11:8] > 6 ? 4'd6 : weighted_sum[265][11:8]);
assign out[266] = (weighted_sum[266][12]==1) ? 4'd0 : (weighted_sum[266][11:8] > 6 ? 4'd6 : weighted_sum[266][11:8]);
assign out[267] = (weighted_sum[267][12]==1) ? 4'd0 : (weighted_sum[267][11:8] > 6 ? 4'd6 : weighted_sum[267][11:8]);
assign out[268] = (weighted_sum[268][12]==1) ? 4'd0 : (weighted_sum[268][11:8] > 6 ? 4'd6 : weighted_sum[268][11:8]);
assign out[269] = (weighted_sum[269][12]==1) ? 4'd0 : (weighted_sum[269][11:8] > 6 ? 4'd6 : weighted_sum[269][11:8]);
assign out[270] = (weighted_sum[270][12]==1) ? 4'd0 : (weighted_sum[270][11:8] > 6 ? 4'd6 : weighted_sum[270][11:8]);
assign out[271] = (weighted_sum[271][12]==1) ? 4'd0 : (weighted_sum[271][11:8] > 6 ? 4'd6 : weighted_sum[271][11:8]);
assign out[272] = (weighted_sum[272][12]==1) ? 4'd0 : (weighted_sum[272][11:8] > 6 ? 4'd6 : weighted_sum[272][11:8]);
assign out[273] = (weighted_sum[273][12]==1) ? 4'd0 : (weighted_sum[273][11:8] > 6 ? 4'd6 : weighted_sum[273][11:8]);
assign out[274] = (weighted_sum[274][12]==1) ? 4'd0 : (weighted_sum[274][11:8] > 6 ? 4'd6 : weighted_sum[274][11:8]);
assign out[275] = (weighted_sum[275][12]==1) ? 4'd0 : (weighted_sum[275][11:8] > 6 ? 4'd6 : weighted_sum[275][11:8]);
assign out[276] = (weighted_sum[276][12]==1) ? 4'd0 : (weighted_sum[276][11:8] > 6 ? 4'd6 : weighted_sum[276][11:8]);
assign out[277] = (weighted_sum[277][12]==1) ? 4'd0 : (weighted_sum[277][11:8] > 6 ? 4'd6 : weighted_sum[277][11:8]);
assign out[278] = (weighted_sum[278][12]==1) ? 4'd0 : (weighted_sum[278][11:8] > 6 ? 4'd6 : weighted_sum[278][11:8]);
assign out[279] = (weighted_sum[279][12]==1) ? 4'd0 : (weighted_sum[279][11:8] > 6 ? 4'd6 : weighted_sum[279][11:8]);
assign out[280] = (weighted_sum[280][12]==1) ? 4'd0 : (weighted_sum[280][11:8] > 6 ? 4'd6 : weighted_sum[280][11:8]);
assign out[281] = (weighted_sum[281][12]==1) ? 4'd0 : (weighted_sum[281][11:8] > 6 ? 4'd6 : weighted_sum[281][11:8]);
assign out[282] = (weighted_sum[282][12]==1) ? 4'd0 : (weighted_sum[282][11:8] > 6 ? 4'd6 : weighted_sum[282][11:8]);
assign out[283] = (weighted_sum[283][12]==1) ? 4'd0 : (weighted_sum[283][11:8] > 6 ? 4'd6 : weighted_sum[283][11:8]);
assign out[284] = (weighted_sum[284][12]==1) ? 4'd0 : (weighted_sum[284][11:8] > 6 ? 4'd6 : weighted_sum[284][11:8]);
assign out[285] = (weighted_sum[285][12]==1) ? 4'd0 : (weighted_sum[285][11:8] > 6 ? 4'd6 : weighted_sum[285][11:8]);
assign out[286] = (weighted_sum[286][12]==1) ? 4'd0 : (weighted_sum[286][11:8] > 6 ? 4'd6 : weighted_sum[286][11:8]);
assign out[287] = (weighted_sum[287][12]==1) ? 4'd0 : (weighted_sum[287][11:8] > 6 ? 4'd6 : weighted_sum[287][11:8]);
assign out[288] = (weighted_sum[288][12]==1) ? 4'd0 : (weighted_sum[288][11:8] > 6 ? 4'd6 : weighted_sum[288][11:8]);
assign out[289] = (weighted_sum[289][12]==1) ? 4'd0 : (weighted_sum[289][11:8] > 6 ? 4'd6 : weighted_sum[289][11:8]);
assign out[290] = (weighted_sum[290][12]==1) ? 4'd0 : (weighted_sum[290][11:8] > 6 ? 4'd6 : weighted_sum[290][11:8]);
assign out[291] = (weighted_sum[291][12]==1) ? 4'd0 : (weighted_sum[291][11:8] > 6 ? 4'd6 : weighted_sum[291][11:8]);
assign out[292] = (weighted_sum[292][12]==1) ? 4'd0 : (weighted_sum[292][11:8] > 6 ? 4'd6 : weighted_sum[292][11:8]);
assign out[293] = (weighted_sum[293][12]==1) ? 4'd0 : (weighted_sum[293][11:8] > 6 ? 4'd6 : weighted_sum[293][11:8]);
assign out[294] = (weighted_sum[294][12]==1) ? 4'd0 : (weighted_sum[294][11:8] > 6 ? 4'd6 : weighted_sum[294][11:8]);
assign out[295] = (weighted_sum[295][12]==1) ? 4'd0 : (weighted_sum[295][11:8] > 6 ? 4'd6 : weighted_sum[295][11:8]);
assign out[296] = (weighted_sum[296][12]==1) ? 4'd0 : (weighted_sum[296][11:8] > 6 ? 4'd6 : weighted_sum[296][11:8]);
assign out[297] = (weighted_sum[297][12]==1) ? 4'd0 : (weighted_sum[297][11:8] > 6 ? 4'd6 : weighted_sum[297][11:8]);
assign out[298] = (weighted_sum[298][12]==1) ? 4'd0 : (weighted_sum[298][11:8] > 6 ? 4'd6 : weighted_sum[298][11:8]);
assign out[299] = (weighted_sum[299][12]==1) ? 4'd0 : (weighted_sum[299][11:8] > 6 ? 4'd6 : weighted_sum[299][11:8]);
assign out[300] = (weighted_sum[300][12]==1) ? 4'd0 : (weighted_sum[300][11:8] > 6 ? 4'd6 : weighted_sum[300][11:8]);
assign out[301] = (weighted_sum[301][12]==1) ? 4'd0 : (weighted_sum[301][11:8] > 6 ? 4'd6 : weighted_sum[301][11:8]);
assign out[302] = (weighted_sum[302][12]==1) ? 4'd0 : (weighted_sum[302][11:8] > 6 ? 4'd6 : weighted_sum[302][11:8]);
assign out[303] = (weighted_sum[303][12]==1) ? 4'd0 : (weighted_sum[303][11:8] > 6 ? 4'd6 : weighted_sum[303][11:8]);
assign out[304] = (weighted_sum[304][12]==1) ? 4'd0 : (weighted_sum[304][11:8] > 6 ? 4'd6 : weighted_sum[304][11:8]);
assign out[305] = (weighted_sum[305][12]==1) ? 4'd0 : (weighted_sum[305][11:8] > 6 ? 4'd6 : weighted_sum[305][11:8]);
assign out[306] = (weighted_sum[306][12]==1) ? 4'd0 : (weighted_sum[306][11:8] > 6 ? 4'd6 : weighted_sum[306][11:8]);
assign out[307] = (weighted_sum[307][12]==1) ? 4'd0 : (weighted_sum[307][11:8] > 6 ? 4'd6 : weighted_sum[307][11:8]);
assign out[308] = (weighted_sum[308][12]==1) ? 4'd0 : (weighted_sum[308][11:8] > 6 ? 4'd6 : weighted_sum[308][11:8]);
assign out[309] = (weighted_sum[309][12]==1) ? 4'd0 : (weighted_sum[309][11:8] > 6 ? 4'd6 : weighted_sum[309][11:8]);
assign out[310] = (weighted_sum[310][12]==1) ? 4'd0 : (weighted_sum[310][11:8] > 6 ? 4'd6 : weighted_sum[310][11:8]);
assign out[311] = (weighted_sum[311][12]==1) ? 4'd0 : (weighted_sum[311][11:8] > 6 ? 4'd6 : weighted_sum[311][11:8]);
assign out[312] = (weighted_sum[312][12]==1) ? 4'd0 : (weighted_sum[312][11:8] > 6 ? 4'd6 : weighted_sum[312][11:8]);
assign out[313] = (weighted_sum[313][12]==1) ? 4'd0 : (weighted_sum[313][11:8] > 6 ? 4'd6 : weighted_sum[313][11:8]);
assign out[314] = (weighted_sum[314][12]==1) ? 4'd0 : (weighted_sum[314][11:8] > 6 ? 4'd6 : weighted_sum[314][11:8]);
assign out[315] = (weighted_sum[315][12]==1) ? 4'd0 : (weighted_sum[315][11:8] > 6 ? 4'd6 : weighted_sum[315][11:8]);
assign out[316] = (weighted_sum[316][12]==1) ? 4'd0 : (weighted_sum[316][11:8] > 6 ? 4'd6 : weighted_sum[316][11:8]);
assign out[317] = (weighted_sum[317][12]==1) ? 4'd0 : (weighted_sum[317][11:8] > 6 ? 4'd6 : weighted_sum[317][11:8]);
assign out[318] = (weighted_sum[318][12]==1) ? 4'd0 : (weighted_sum[318][11:8] > 6 ? 4'd6 : weighted_sum[318][11:8]);
assign out[319] = (weighted_sum[319][12]==1) ? 4'd0 : (weighted_sum[319][11:8] > 6 ? 4'd6 : weighted_sum[319][11:8]);
assign out[320] = (weighted_sum[320][12]==1) ? 4'd0 : (weighted_sum[320][11:8] > 6 ? 4'd6 : weighted_sum[320][11:8]);
assign out[321] = (weighted_sum[321][12]==1) ? 4'd0 : (weighted_sum[321][11:8] > 6 ? 4'd6 : weighted_sum[321][11:8]);
assign out[322] = (weighted_sum[322][12]==1) ? 4'd0 : (weighted_sum[322][11:8] > 6 ? 4'd6 : weighted_sum[322][11:8]);
assign out[323] = (weighted_sum[323][12]==1) ? 4'd0 : (weighted_sum[323][11:8] > 6 ? 4'd6 : weighted_sum[323][11:8]);
assign out[324] = (weighted_sum[324][12]==1) ? 4'd0 : (weighted_sum[324][11:8] > 6 ? 4'd6 : weighted_sum[324][11:8]);
assign out[325] = (weighted_sum[325][12]==1) ? 4'd0 : (weighted_sum[325][11:8] > 6 ? 4'd6 : weighted_sum[325][11:8]);
assign out[326] = (weighted_sum[326][12]==1) ? 4'd0 : (weighted_sum[326][11:8] > 6 ? 4'd6 : weighted_sum[326][11:8]);
assign out[327] = (weighted_sum[327][12]==1) ? 4'd0 : (weighted_sum[327][11:8] > 6 ? 4'd6 : weighted_sum[327][11:8]);
assign out[328] = (weighted_sum[328][12]==1) ? 4'd0 : (weighted_sum[328][11:8] > 6 ? 4'd6 : weighted_sum[328][11:8]);
assign out[329] = (weighted_sum[329][12]==1) ? 4'd0 : (weighted_sum[329][11:8] > 6 ? 4'd6 : weighted_sum[329][11:8]);
assign out[330] = (weighted_sum[330][12]==1) ? 4'd0 : (weighted_sum[330][11:8] > 6 ? 4'd6 : weighted_sum[330][11:8]);
assign out[331] = (weighted_sum[331][12]==1) ? 4'd0 : (weighted_sum[331][11:8] > 6 ? 4'd6 : weighted_sum[331][11:8]);
assign out[332] = (weighted_sum[332][12]==1) ? 4'd0 : (weighted_sum[332][11:8] > 6 ? 4'd6 : weighted_sum[332][11:8]);
assign out[333] = (weighted_sum[333][12]==1) ? 4'd0 : (weighted_sum[333][11:8] > 6 ? 4'd6 : weighted_sum[333][11:8]);
assign out[334] = (weighted_sum[334][12]==1) ? 4'd0 : (weighted_sum[334][11:8] > 6 ? 4'd6 : weighted_sum[334][11:8]);
assign out[335] = (weighted_sum[335][12]==1) ? 4'd0 : (weighted_sum[335][11:8] > 6 ? 4'd6 : weighted_sum[335][11:8]);
assign out[336] = (weighted_sum[336][12]==1) ? 4'd0 : (weighted_sum[336][11:8] > 6 ? 4'd6 : weighted_sum[336][11:8]);
assign out[337] = (weighted_sum[337][12]==1) ? 4'd0 : (weighted_sum[337][11:8] > 6 ? 4'd6 : weighted_sum[337][11:8]);
assign out[338] = (weighted_sum[338][12]==1) ? 4'd0 : (weighted_sum[338][11:8] > 6 ? 4'd6 : weighted_sum[338][11:8]);
assign out[339] = (weighted_sum[339][12]==1) ? 4'd0 : (weighted_sum[339][11:8] > 6 ? 4'd6 : weighted_sum[339][11:8]);
assign out[340] = (weighted_sum[340][12]==1) ? 4'd0 : (weighted_sum[340][11:8] > 6 ? 4'd6 : weighted_sum[340][11:8]);
assign out[341] = (weighted_sum[341][12]==1) ? 4'd0 : (weighted_sum[341][11:8] > 6 ? 4'd6 : weighted_sum[341][11:8]);
assign out[342] = (weighted_sum[342][12]==1) ? 4'd0 : (weighted_sum[342][11:8] > 6 ? 4'd6 : weighted_sum[342][11:8]);
assign out[343] = (weighted_sum[343][12]==1) ? 4'd0 : (weighted_sum[343][11:8] > 6 ? 4'd6 : weighted_sum[343][11:8]);
assign out[344] = (weighted_sum[344][12]==1) ? 4'd0 : (weighted_sum[344][11:8] > 6 ? 4'd6 : weighted_sum[344][11:8]);
assign out[345] = (weighted_sum[345][12]==1) ? 4'd0 : (weighted_sum[345][11:8] > 6 ? 4'd6 : weighted_sum[345][11:8]);
assign out[346] = (weighted_sum[346][12]==1) ? 4'd0 : (weighted_sum[346][11:8] > 6 ? 4'd6 : weighted_sum[346][11:8]);
assign out[347] = (weighted_sum[347][12]==1) ? 4'd0 : (weighted_sum[347][11:8] > 6 ? 4'd6 : weighted_sum[347][11:8]);
assign out[348] = (weighted_sum[348][12]==1) ? 4'd0 : (weighted_sum[348][11:8] > 6 ? 4'd6 : weighted_sum[348][11:8]);
assign out[349] = (weighted_sum[349][12]==1) ? 4'd0 : (weighted_sum[349][11:8] > 6 ? 4'd6 : weighted_sum[349][11:8]);
assign out[350] = (weighted_sum[350][12]==1) ? 4'd0 : (weighted_sum[350][11:8] > 6 ? 4'd6 : weighted_sum[350][11:8]);
assign out[351] = (weighted_sum[351][12]==1) ? 4'd0 : (weighted_sum[351][11:8] > 6 ? 4'd6 : weighted_sum[351][11:8]);
assign out[352] = (weighted_sum[352][12]==1) ? 4'd0 : (weighted_sum[352][11:8] > 6 ? 4'd6 : weighted_sum[352][11:8]);
assign out[353] = (weighted_sum[353][12]==1) ? 4'd0 : (weighted_sum[353][11:8] > 6 ? 4'd6 : weighted_sum[353][11:8]);
assign out[354] = (weighted_sum[354][12]==1) ? 4'd0 : (weighted_sum[354][11:8] > 6 ? 4'd6 : weighted_sum[354][11:8]);
assign out[355] = (weighted_sum[355][12]==1) ? 4'd0 : (weighted_sum[355][11:8] > 6 ? 4'd6 : weighted_sum[355][11:8]);
assign out[356] = (weighted_sum[356][12]==1) ? 4'd0 : (weighted_sum[356][11:8] > 6 ? 4'd6 : weighted_sum[356][11:8]);
assign out[357] = (weighted_sum[357][12]==1) ? 4'd0 : (weighted_sum[357][11:8] > 6 ? 4'd6 : weighted_sum[357][11:8]);
assign out[358] = (weighted_sum[358][12]==1) ? 4'd0 : (weighted_sum[358][11:8] > 6 ? 4'd6 : weighted_sum[358][11:8]);
assign out[359] = (weighted_sum[359][12]==1) ? 4'd0 : (weighted_sum[359][11:8] > 6 ? 4'd6 : weighted_sum[359][11:8]);
assign out[360] = (weighted_sum[360][12]==1) ? 4'd0 : (weighted_sum[360][11:8] > 6 ? 4'd6 : weighted_sum[360][11:8]);
assign out[361] = (weighted_sum[361][12]==1) ? 4'd0 : (weighted_sum[361][11:8] > 6 ? 4'd6 : weighted_sum[361][11:8]);
assign out[362] = (weighted_sum[362][12]==1) ? 4'd0 : (weighted_sum[362][11:8] > 6 ? 4'd6 : weighted_sum[362][11:8]);
assign out[363] = (weighted_sum[363][12]==1) ? 4'd0 : (weighted_sum[363][11:8] > 6 ? 4'd6 : weighted_sum[363][11:8]);
assign out[364] = (weighted_sum[364][12]==1) ? 4'd0 : (weighted_sum[364][11:8] > 6 ? 4'd6 : weighted_sum[364][11:8]);
assign out[365] = (weighted_sum[365][12]==1) ? 4'd0 : (weighted_sum[365][11:8] > 6 ? 4'd6 : weighted_sum[365][11:8]);
assign out[366] = (weighted_sum[366][12]==1) ? 4'd0 : (weighted_sum[366][11:8] > 6 ? 4'd6 : weighted_sum[366][11:8]);
assign out[367] = (weighted_sum[367][12]==1) ? 4'd0 : (weighted_sum[367][11:8] > 6 ? 4'd6 : weighted_sum[367][11:8]);
assign out[368] = (weighted_sum[368][12]==1) ? 4'd0 : (weighted_sum[368][11:8] > 6 ? 4'd6 : weighted_sum[368][11:8]);
assign out[369] = (weighted_sum[369][12]==1) ? 4'd0 : (weighted_sum[369][11:8] > 6 ? 4'd6 : weighted_sum[369][11:8]);
assign out[370] = (weighted_sum[370][12]==1) ? 4'd0 : (weighted_sum[370][11:8] > 6 ? 4'd6 : weighted_sum[370][11:8]);
assign out[371] = (weighted_sum[371][12]==1) ? 4'd0 : (weighted_sum[371][11:8] > 6 ? 4'd6 : weighted_sum[371][11:8]);
assign out[372] = (weighted_sum[372][12]==1) ? 4'd0 : (weighted_sum[372][11:8] > 6 ? 4'd6 : weighted_sum[372][11:8]);
assign out[373] = (weighted_sum[373][12]==1) ? 4'd0 : (weighted_sum[373][11:8] > 6 ? 4'd6 : weighted_sum[373][11:8]);
assign out[374] = (weighted_sum[374][12]==1) ? 4'd0 : (weighted_sum[374][11:8] > 6 ? 4'd6 : weighted_sum[374][11:8]);
assign out[375] = (weighted_sum[375][12]==1) ? 4'd0 : (weighted_sum[375][11:8] > 6 ? 4'd6 : weighted_sum[375][11:8]);
assign out[376] = (weighted_sum[376][12]==1) ? 4'd0 : (weighted_sum[376][11:8] > 6 ? 4'd6 : weighted_sum[376][11:8]);
assign out[377] = (weighted_sum[377][12]==1) ? 4'd0 : (weighted_sum[377][11:8] > 6 ? 4'd6 : weighted_sum[377][11:8]);
assign out[378] = (weighted_sum[378][12]==1) ? 4'd0 : (weighted_sum[378][11:8] > 6 ? 4'd6 : weighted_sum[378][11:8]);
assign out[379] = (weighted_sum[379][12]==1) ? 4'd0 : (weighted_sum[379][11:8] > 6 ? 4'd6 : weighted_sum[379][11:8]);
assign out[380] = (weighted_sum[380][12]==1) ? 4'd0 : (weighted_sum[380][11:8] > 6 ? 4'd6 : weighted_sum[380][11:8]);
assign out[381] = (weighted_sum[381][12]==1) ? 4'd0 : (weighted_sum[381][11:8] > 6 ? 4'd6 : weighted_sum[381][11:8]);
assign out[382] = (weighted_sum[382][12]==1) ? 4'd0 : (weighted_sum[382][11:8] > 6 ? 4'd6 : weighted_sum[382][11:8]);
assign out[383] = (weighted_sum[383][12]==1) ? 4'd0 : (weighted_sum[383][11:8] > 6 ? 4'd6 : weighted_sum[383][11:8]);
assign out[384] = (weighted_sum[384][12]==1) ? 4'd0 : (weighted_sum[384][11:8] > 6 ? 4'd6 : weighted_sum[384][11:8]);
assign out[385] = (weighted_sum[385][12]==1) ? 4'd0 : (weighted_sum[385][11:8] > 6 ? 4'd6 : weighted_sum[385][11:8]);
assign out[386] = (weighted_sum[386][12]==1) ? 4'd0 : (weighted_sum[386][11:8] > 6 ? 4'd6 : weighted_sum[386][11:8]);
assign out[387] = (weighted_sum[387][12]==1) ? 4'd0 : (weighted_sum[387][11:8] > 6 ? 4'd6 : weighted_sum[387][11:8]);
assign out[388] = (weighted_sum[388][12]==1) ? 4'd0 : (weighted_sum[388][11:8] > 6 ? 4'd6 : weighted_sum[388][11:8]);
assign out[389] = (weighted_sum[389][12]==1) ? 4'd0 : (weighted_sum[389][11:8] > 6 ? 4'd6 : weighted_sum[389][11:8]);
assign out[390] = (weighted_sum[390][12]==1) ? 4'd0 : (weighted_sum[390][11:8] > 6 ? 4'd6 : weighted_sum[390][11:8]);
assign out[391] = (weighted_sum[391][12]==1) ? 4'd0 : (weighted_sum[391][11:8] > 6 ? 4'd6 : weighted_sum[391][11:8]);
assign out[392] = (weighted_sum[392][12]==1) ? 4'd0 : (weighted_sum[392][11:8] > 6 ? 4'd6 : weighted_sum[392][11:8]);
assign out[393] = (weighted_sum[393][12]==1) ? 4'd0 : (weighted_sum[393][11:8] > 6 ? 4'd6 : weighted_sum[393][11:8]);
assign out[394] = (weighted_sum[394][12]==1) ? 4'd0 : (weighted_sum[394][11:8] > 6 ? 4'd6 : weighted_sum[394][11:8]);
assign out[395] = (weighted_sum[395][12]==1) ? 4'd0 : (weighted_sum[395][11:8] > 6 ? 4'd6 : weighted_sum[395][11:8]);
assign out[396] = (weighted_sum[396][12]==1) ? 4'd0 : (weighted_sum[396][11:8] > 6 ? 4'd6 : weighted_sum[396][11:8]);
assign out[397] = (weighted_sum[397][12]==1) ? 4'd0 : (weighted_sum[397][11:8] > 6 ? 4'd6 : weighted_sum[397][11:8]);
assign out[398] = (weighted_sum[398][12]==1) ? 4'd0 : (weighted_sum[398][11:8] > 6 ? 4'd6 : weighted_sum[398][11:8]);
assign out[399] = (weighted_sum[399][12]==1) ? 4'd0 : (weighted_sum[399][11:8] > 6 ? 4'd6 : weighted_sum[399][11:8]);
assign out[400] = (weighted_sum[400][12]==1) ? 4'd0 : (weighted_sum[400][11:8] > 6 ? 4'd6 : weighted_sum[400][11:8]);
assign out[401] = (weighted_sum[401][12]==1) ? 4'd0 : (weighted_sum[401][11:8] > 6 ? 4'd6 : weighted_sum[401][11:8]);
assign out[402] = (weighted_sum[402][12]==1) ? 4'd0 : (weighted_sum[402][11:8] > 6 ? 4'd6 : weighted_sum[402][11:8]);
assign out[403] = (weighted_sum[403][12]==1) ? 4'd0 : (weighted_sum[403][11:8] > 6 ? 4'd6 : weighted_sum[403][11:8]);
assign out[404] = (weighted_sum[404][12]==1) ? 4'd0 : (weighted_sum[404][11:8] > 6 ? 4'd6 : weighted_sum[404][11:8]);
assign out[405] = (weighted_sum[405][12]==1) ? 4'd0 : (weighted_sum[405][11:8] > 6 ? 4'd6 : weighted_sum[405][11:8]);
assign out[406] = (weighted_sum[406][12]==1) ? 4'd0 : (weighted_sum[406][11:8] > 6 ? 4'd6 : weighted_sum[406][11:8]);
assign out[407] = (weighted_sum[407][12]==1) ? 4'd0 : (weighted_sum[407][11:8] > 6 ? 4'd6 : weighted_sum[407][11:8]);
assign out[408] = (weighted_sum[408][12]==1) ? 4'd0 : (weighted_sum[408][11:8] > 6 ? 4'd6 : weighted_sum[408][11:8]);
assign out[409] = (weighted_sum[409][12]==1) ? 4'd0 : (weighted_sum[409][11:8] > 6 ? 4'd6 : weighted_sum[409][11:8]);
assign out[410] = (weighted_sum[410][12]==1) ? 4'd0 : (weighted_sum[410][11:8] > 6 ? 4'd6 : weighted_sum[410][11:8]);
assign out[411] = (weighted_sum[411][12]==1) ? 4'd0 : (weighted_sum[411][11:8] > 6 ? 4'd6 : weighted_sum[411][11:8]);
assign out[412] = (weighted_sum[412][12]==1) ? 4'd0 : (weighted_sum[412][11:8] > 6 ? 4'd6 : weighted_sum[412][11:8]);
assign out[413] = (weighted_sum[413][12]==1) ? 4'd0 : (weighted_sum[413][11:8] > 6 ? 4'd6 : weighted_sum[413][11:8]);
assign out[414] = (weighted_sum[414][12]==1) ? 4'd0 : (weighted_sum[414][11:8] > 6 ? 4'd6 : weighted_sum[414][11:8]);
assign out[415] = (weighted_sum[415][12]==1) ? 4'd0 : (weighted_sum[415][11:8] > 6 ? 4'd6 : weighted_sum[415][11:8]);
assign out[416] = (weighted_sum[416][12]==1) ? 4'd0 : (weighted_sum[416][11:8] > 6 ? 4'd6 : weighted_sum[416][11:8]);
assign out[417] = (weighted_sum[417][12]==1) ? 4'd0 : (weighted_sum[417][11:8] > 6 ? 4'd6 : weighted_sum[417][11:8]);
assign out[418] = (weighted_sum[418][12]==1) ? 4'd0 : (weighted_sum[418][11:8] > 6 ? 4'd6 : weighted_sum[418][11:8]);
assign out[419] = (weighted_sum[419][12]==1) ? 4'd0 : (weighted_sum[419][11:8] > 6 ? 4'd6 : weighted_sum[419][11:8]);
assign out[420] = (weighted_sum[420][12]==1) ? 4'd0 : (weighted_sum[420][11:8] > 6 ? 4'd6 : weighted_sum[420][11:8]);
assign out[421] = (weighted_sum[421][12]==1) ? 4'd0 : (weighted_sum[421][11:8] > 6 ? 4'd6 : weighted_sum[421][11:8]);
assign out[422] = (weighted_sum[422][12]==1) ? 4'd0 : (weighted_sum[422][11:8] > 6 ? 4'd6 : weighted_sum[422][11:8]);
assign out[423] = (weighted_sum[423][12]==1) ? 4'd0 : (weighted_sum[423][11:8] > 6 ? 4'd6 : weighted_sum[423][11:8]);
assign out[424] = (weighted_sum[424][12]==1) ? 4'd0 : (weighted_sum[424][11:8] > 6 ? 4'd6 : weighted_sum[424][11:8]);
assign out[425] = (weighted_sum[425][12]==1) ? 4'd0 : (weighted_sum[425][11:8] > 6 ? 4'd6 : weighted_sum[425][11:8]);
assign out[426] = (weighted_sum[426][12]==1) ? 4'd0 : (weighted_sum[426][11:8] > 6 ? 4'd6 : weighted_sum[426][11:8]);
assign out[427] = (weighted_sum[427][12]==1) ? 4'd0 : (weighted_sum[427][11:8] > 6 ? 4'd6 : weighted_sum[427][11:8]);
assign out[428] = (weighted_sum[428][12]==1) ? 4'd0 : (weighted_sum[428][11:8] > 6 ? 4'd6 : weighted_sum[428][11:8]);
assign out[429] = (weighted_sum[429][12]==1) ? 4'd0 : (weighted_sum[429][11:8] > 6 ? 4'd6 : weighted_sum[429][11:8]);
assign out[430] = (weighted_sum[430][12]==1) ? 4'd0 : (weighted_sum[430][11:8] > 6 ? 4'd6 : weighted_sum[430][11:8]);
assign out[431] = (weighted_sum[431][12]==1) ? 4'd0 : (weighted_sum[431][11:8] > 6 ? 4'd6 : weighted_sum[431][11:8]);
assign out[432] = (weighted_sum[432][12]==1) ? 4'd0 : (weighted_sum[432][11:8] > 6 ? 4'd6 : weighted_sum[432][11:8]);
assign out[433] = (weighted_sum[433][12]==1) ? 4'd0 : (weighted_sum[433][11:8] > 6 ? 4'd6 : weighted_sum[433][11:8]);
assign out[434] = (weighted_sum[434][12]==1) ? 4'd0 : (weighted_sum[434][11:8] > 6 ? 4'd6 : weighted_sum[434][11:8]);
assign out[435] = (weighted_sum[435][12]==1) ? 4'd0 : (weighted_sum[435][11:8] > 6 ? 4'd6 : weighted_sum[435][11:8]);
assign out[436] = (weighted_sum[436][12]==1) ? 4'd0 : (weighted_sum[436][11:8] > 6 ? 4'd6 : weighted_sum[436][11:8]);
assign out[437] = (weighted_sum[437][12]==1) ? 4'd0 : (weighted_sum[437][11:8] > 6 ? 4'd6 : weighted_sum[437][11:8]);
assign out[438] = (weighted_sum[438][12]==1) ? 4'd0 : (weighted_sum[438][11:8] > 6 ? 4'd6 : weighted_sum[438][11:8]);
assign out[439] = (weighted_sum[439][12]==1) ? 4'd0 : (weighted_sum[439][11:8] > 6 ? 4'd6 : weighted_sum[439][11:8]);
assign out[440] = (weighted_sum[440][12]==1) ? 4'd0 : (weighted_sum[440][11:8] > 6 ? 4'd6 : weighted_sum[440][11:8]);
assign out[441] = (weighted_sum[441][12]==1) ? 4'd0 : (weighted_sum[441][11:8] > 6 ? 4'd6 : weighted_sum[441][11:8]);
assign out[442] = (weighted_sum[442][12]==1) ? 4'd0 : (weighted_sum[442][11:8] > 6 ? 4'd6 : weighted_sum[442][11:8]);
assign out[443] = (weighted_sum[443][12]==1) ? 4'd0 : (weighted_sum[443][11:8] > 6 ? 4'd6 : weighted_sum[443][11:8]);
assign out[444] = (weighted_sum[444][12]==1) ? 4'd0 : (weighted_sum[444][11:8] > 6 ? 4'd6 : weighted_sum[444][11:8]);
assign out[445] = (weighted_sum[445][12]==1) ? 4'd0 : (weighted_sum[445][11:8] > 6 ? 4'd6 : weighted_sum[445][11:8]);
assign out[446] = (weighted_sum[446][12]==1) ? 4'd0 : (weighted_sum[446][11:8] > 6 ? 4'd6 : weighted_sum[446][11:8]);
assign out[447] = (weighted_sum[447][12]==1) ? 4'd0 : (weighted_sum[447][11:8] > 6 ? 4'd6 : weighted_sum[447][11:8]);
assign out[448] = (weighted_sum[448][12]==1) ? 4'd0 : (weighted_sum[448][11:8] > 6 ? 4'd6 : weighted_sum[448][11:8]);
assign out[449] = (weighted_sum[449][12]==1) ? 4'd0 : (weighted_sum[449][11:8] > 6 ? 4'd6 : weighted_sum[449][11:8]);
assign out[450] = (weighted_sum[450][12]==1) ? 4'd0 : (weighted_sum[450][11:8] > 6 ? 4'd6 : weighted_sum[450][11:8]);
assign out[451] = (weighted_sum[451][12]==1) ? 4'd0 : (weighted_sum[451][11:8] > 6 ? 4'd6 : weighted_sum[451][11:8]);
assign out[452] = (weighted_sum[452][12]==1) ? 4'd0 : (weighted_sum[452][11:8] > 6 ? 4'd6 : weighted_sum[452][11:8]);
assign out[453] = (weighted_sum[453][12]==1) ? 4'd0 : (weighted_sum[453][11:8] > 6 ? 4'd6 : weighted_sum[453][11:8]);
assign out[454] = (weighted_sum[454][12]==1) ? 4'd0 : (weighted_sum[454][11:8] > 6 ? 4'd6 : weighted_sum[454][11:8]);
assign out[455] = (weighted_sum[455][12]==1) ? 4'd0 : (weighted_sum[455][11:8] > 6 ? 4'd6 : weighted_sum[455][11:8]);
assign out[456] = (weighted_sum[456][12]==1) ? 4'd0 : (weighted_sum[456][11:8] > 6 ? 4'd6 : weighted_sum[456][11:8]);
assign out[457] = (weighted_sum[457][12]==1) ? 4'd0 : (weighted_sum[457][11:8] > 6 ? 4'd6 : weighted_sum[457][11:8]);
assign out[458] = (weighted_sum[458][12]==1) ? 4'd0 : (weighted_sum[458][11:8] > 6 ? 4'd6 : weighted_sum[458][11:8]);
assign out[459] = (weighted_sum[459][12]==1) ? 4'd0 : (weighted_sum[459][11:8] > 6 ? 4'd6 : weighted_sum[459][11:8]);
assign out[460] = (weighted_sum[460][12]==1) ? 4'd0 : (weighted_sum[460][11:8] > 6 ? 4'd6 : weighted_sum[460][11:8]);
assign out[461] = (weighted_sum[461][12]==1) ? 4'd0 : (weighted_sum[461][11:8] > 6 ? 4'd6 : weighted_sum[461][11:8]);
assign out[462] = (weighted_sum[462][12]==1) ? 4'd0 : (weighted_sum[462][11:8] > 6 ? 4'd6 : weighted_sum[462][11:8]);
assign out[463] = (weighted_sum[463][12]==1) ? 4'd0 : (weighted_sum[463][11:8] > 6 ? 4'd6 : weighted_sum[463][11:8]);
assign out[464] = (weighted_sum[464][12]==1) ? 4'd0 : (weighted_sum[464][11:8] > 6 ? 4'd6 : weighted_sum[464][11:8]);
assign out[465] = (weighted_sum[465][12]==1) ? 4'd0 : (weighted_sum[465][11:8] > 6 ? 4'd6 : weighted_sum[465][11:8]);
assign out[466] = (weighted_sum[466][12]==1) ? 4'd0 : (weighted_sum[466][11:8] > 6 ? 4'd6 : weighted_sum[466][11:8]);
assign out[467] = (weighted_sum[467][12]==1) ? 4'd0 : (weighted_sum[467][11:8] > 6 ? 4'd6 : weighted_sum[467][11:8]);
assign out[468] = (weighted_sum[468][12]==1) ? 4'd0 : (weighted_sum[468][11:8] > 6 ? 4'd6 : weighted_sum[468][11:8]);
assign out[469] = (weighted_sum[469][12]==1) ? 4'd0 : (weighted_sum[469][11:8] > 6 ? 4'd6 : weighted_sum[469][11:8]);
assign out[470] = (weighted_sum[470][12]==1) ? 4'd0 : (weighted_sum[470][11:8] > 6 ? 4'd6 : weighted_sum[470][11:8]);
assign out[471] = (weighted_sum[471][12]==1) ? 4'd0 : (weighted_sum[471][11:8] > 6 ? 4'd6 : weighted_sum[471][11:8]);
assign out[472] = (weighted_sum[472][12]==1) ? 4'd0 : (weighted_sum[472][11:8] > 6 ? 4'd6 : weighted_sum[472][11:8]);
assign out[473] = (weighted_sum[473][12]==1) ? 4'd0 : (weighted_sum[473][11:8] > 6 ? 4'd6 : weighted_sum[473][11:8]);
assign out[474] = (weighted_sum[474][12]==1) ? 4'd0 : (weighted_sum[474][11:8] > 6 ? 4'd6 : weighted_sum[474][11:8]);
assign out[475] = (weighted_sum[475][12]==1) ? 4'd0 : (weighted_sum[475][11:8] > 6 ? 4'd6 : weighted_sum[475][11:8]);
assign out[476] = (weighted_sum[476][12]==1) ? 4'd0 : (weighted_sum[476][11:8] > 6 ? 4'd6 : weighted_sum[476][11:8]);
assign out[477] = (weighted_sum[477][12]==1) ? 4'd0 : (weighted_sum[477][11:8] > 6 ? 4'd6 : weighted_sum[477][11:8]);
assign out[478] = (weighted_sum[478][12]==1) ? 4'd0 : (weighted_sum[478][11:8] > 6 ? 4'd6 : weighted_sum[478][11:8]);
assign out[479] = (weighted_sum[479][12]==1) ? 4'd0 : (weighted_sum[479][11:8] > 6 ? 4'd6 : weighted_sum[479][11:8]);
assign out[480] = (weighted_sum[480][12]==1) ? 4'd0 : (weighted_sum[480][11:8] > 6 ? 4'd6 : weighted_sum[480][11:8]);
assign out[481] = (weighted_sum[481][12]==1) ? 4'd0 : (weighted_sum[481][11:8] > 6 ? 4'd6 : weighted_sum[481][11:8]);
assign out[482] = (weighted_sum[482][12]==1) ? 4'd0 : (weighted_sum[482][11:8] > 6 ? 4'd6 : weighted_sum[482][11:8]);
assign out[483] = (weighted_sum[483][12]==1) ? 4'd0 : (weighted_sum[483][11:8] > 6 ? 4'd6 : weighted_sum[483][11:8]);
assign out[484] = (weighted_sum[484][12]==1) ? 4'd0 : (weighted_sum[484][11:8] > 6 ? 4'd6 : weighted_sum[484][11:8]);
assign out[485] = (weighted_sum[485][12]==1) ? 4'd0 : (weighted_sum[485][11:8] > 6 ? 4'd6 : weighted_sum[485][11:8]);
assign out[486] = (weighted_sum[486][12]==1) ? 4'd0 : (weighted_sum[486][11:8] > 6 ? 4'd6 : weighted_sum[486][11:8]);
assign out[487] = (weighted_sum[487][12]==1) ? 4'd0 : (weighted_sum[487][11:8] > 6 ? 4'd6 : weighted_sum[487][11:8]);
assign out[488] = (weighted_sum[488][12]==1) ? 4'd0 : (weighted_sum[488][11:8] > 6 ? 4'd6 : weighted_sum[488][11:8]);
assign out[489] = (weighted_sum[489][12]==1) ? 4'd0 : (weighted_sum[489][11:8] > 6 ? 4'd6 : weighted_sum[489][11:8]);
assign out[490] = (weighted_sum[490][12]==1) ? 4'd0 : (weighted_sum[490][11:8] > 6 ? 4'd6 : weighted_sum[490][11:8]);
assign out[491] = (weighted_sum[491][12]==1) ? 4'd0 : (weighted_sum[491][11:8] > 6 ? 4'd6 : weighted_sum[491][11:8]);
assign out[492] = (weighted_sum[492][12]==1) ? 4'd0 : (weighted_sum[492][11:8] > 6 ? 4'd6 : weighted_sum[492][11:8]);
assign out[493] = (weighted_sum[493][12]==1) ? 4'd0 : (weighted_sum[493][11:8] > 6 ? 4'd6 : weighted_sum[493][11:8]);
assign out[494] = (weighted_sum[494][12]==1) ? 4'd0 : (weighted_sum[494][11:8] > 6 ? 4'd6 : weighted_sum[494][11:8]);
assign out[495] = (weighted_sum[495][12]==1) ? 4'd0 : (weighted_sum[495][11:8] > 6 ? 4'd6 : weighted_sum[495][11:8]);
assign out[496] = (weighted_sum[496][12]==1) ? 4'd0 : (weighted_sum[496][11:8] > 6 ? 4'd6 : weighted_sum[496][11:8]);
assign out[497] = (weighted_sum[497][12]==1) ? 4'd0 : (weighted_sum[497][11:8] > 6 ? 4'd6 : weighted_sum[497][11:8]);
assign out[498] = (weighted_sum[498][12]==1) ? 4'd0 : (weighted_sum[498][11:8] > 6 ? 4'd6 : weighted_sum[498][11:8]);
assign out[499] = (weighted_sum[499][12]==1) ? 4'd0 : (weighted_sum[499][11:8] > 6 ? 4'd6 : weighted_sum[499][11:8]);
assign out[500] = (weighted_sum[500][12]==1) ? 4'd0 : (weighted_sum[500][11:8] > 6 ? 4'd6 : weighted_sum[500][11:8]);
assign out[501] = (weighted_sum[501][12]==1) ? 4'd0 : (weighted_sum[501][11:8] > 6 ? 4'd6 : weighted_sum[501][11:8]);
assign out[502] = (weighted_sum[502][12]==1) ? 4'd0 : (weighted_sum[502][11:8] > 6 ? 4'd6 : weighted_sum[502][11:8]);
assign out[503] = (weighted_sum[503][12]==1) ? 4'd0 : (weighted_sum[503][11:8] > 6 ? 4'd6 : weighted_sum[503][11:8]);
assign out[504] = (weighted_sum[504][12]==1) ? 4'd0 : (weighted_sum[504][11:8] > 6 ? 4'd6 : weighted_sum[504][11:8]);
assign out[505] = (weighted_sum[505][12]==1) ? 4'd0 : (weighted_sum[505][11:8] > 6 ? 4'd6 : weighted_sum[505][11:8]);
assign out[506] = (weighted_sum[506][12]==1) ? 4'd0 : (weighted_sum[506][11:8] > 6 ? 4'd6 : weighted_sum[506][11:8]);

always_ff @ (posedge clk or posedge rst) begin
	if (rst) begin
		sharing0_r <= 0;
		sharing1_r <= 0;
		sharing2_r <= 0;
		sharing3_r <= 0;
		sharing4_r <= 0;
		sharing5_r <= 0;
		sharing6_r <= 0;
		sharing7_r <= 0;
		sharing8_r <= 0;
		sharing9_r <= 0;
		sharing10_r <= 0;
		sharing11_r <= 0;
		sharing12_r <= 0;
		sharing13_r <= 0;
		sharing14_r <= 0;
		sharing15_r <= 0;
		sharing16_r <= 0;
		sharing17_r <= 0;
		sharing18_r <= 0;
		sharing19_r <= 0;
		sharing20_r <= 0;
		sharing21_r <= 0;
		sharing22_r <= 0;
		sharing23_r <= 0;
		sharing24_r <= 0;
		sharing25_r <= 0;
		sharing26_r <= 0;
		sharing27_r <= 0;
		sharing28_r <= 0;
		sharing29_r <= 0;
		sharing30_r <= 0;
		sharing31_r <= 0;
		sharing32_r <= 0;
		sharing33_r <= 0;
		sharing34_r <= 0;
		sharing35_r <= 0;
		sharing36_r <= 0;
		sharing37_r <= 0;
		sharing38_r <= 0;
		sharing39_r <= 0;
		sharing40_r <= 0;
		sharing41_r <= 0;
		sharing42_r <= 0;
		sharing43_r <= 0;
		sharing44_r <= 0;
		sharing45_r <= 0;
		sharing46_r <= 0;
		sharing47_r <= 0;
		sharing48_r <= 0;
		sharing49_r <= 0;
		sharing50_r <= 0;
		sharing51_r <= 0;
		sharing52_r <= 0;
		sharing53_r <= 0;
		sharing54_r <= 0;
		sharing55_r <= 0;
		sharing56_r <= 0;
		sharing57_r <= 0;
		sharing58_r <= 0;
		sharing59_r <= 0;
		sharing60_r <= 0;
		sharing61_r <= 0;
		sharing62_r <= 0;
		sharing63_r <= 0;
		sharing64_r <= 0;
		sharing65_r <= 0;
		sharing66_r <= 0;
		sharing67_r <= 0;
		sharing68_r <= 0;
		sharing69_r <= 0;
		sharing70_r <= 0;
		sharing71_r <= 0;
		sharing72_r <= 0;
		sharing73_r <= 0;
		sharing74_r <= 0;
		sharing75_r <= 0;
		sharing76_r <= 0;
		sharing77_r <= 0;
		sharing78_r <= 0;
		sharing79_r <= 0;
		sharing80_r <= 0;
		sharing81_r <= 0;
		sharing82_r <= 0;
		sharing83_r <= 0;
		sharing84_r <= 0;
		sharing85_r <= 0;
		sharing86_r <= 0;
		sharing87_r <= 0;
		sharing88_r <= 0;
		sharing89_r <= 0;
		sharing90_r <= 0;
		sharing91_r <= 0;
		sharing92_r <= 0;
		sharing93_r <= 0;
		sharing94_r <= 0;
		sharing95_r <= 0;
		sharing96_r <= 0;
		sharing97_r <= 0;
		sharing98_r <= 0;
		sharing99_r <= 0;
		sharing100_r <= 0;
		sharing101_r <= 0;
		sharing102_r <= 0;
		sharing103_r <= 0;
		sharing104_r <= 0;
		sharing105_r <= 0;
		sharing106_r <= 0;
		sharing107_r <= 0;
		sharing108_r <= 0;
		sharing109_r <= 0;
		sharing110_r <= 0;
		sharing111_r <= 0;
		sharing112_r <= 0;
		sharing113_r <= 0;
		sharing114_r <= 0;
		sharing115_r <= 0;
		sharing116_r <= 0;
		sharing117_r <= 0;
		sharing118_r <= 0;
		sharing119_r <= 0;
		sharing120_r <= 0;
		sharing121_r <= 0;
		sharing122_r <= 0;
		sharing123_r <= 0;
		sharing124_r <= 0;
		sharing125_r <= 0;
		sharing126_r <= 0;
		sharing127_r <= 0;
		sharing128_r <= 0;
		sharing129_r <= 0;
		sharing130_r <= 0;
		sharing131_r <= 0;
		sharing132_r <= 0;
		sharing133_r <= 0;
		sharing134_r <= 0;
		sharing135_r <= 0;
		sharing136_r <= 0;
		sharing137_r <= 0;
		sharing138_r <= 0;
		sharing139_r <= 0;
		sharing140_r <= 0;
		sharing141_r <= 0;
		sharing142_r <= 0;
		sharing143_r <= 0;
		sharing144_r <= 0;
		sharing145_r <= 0;
		sharing146_r <= 0;
		sharing147_r <= 0;
		sharing148_r <= 0;
		sharing149_r <= 0;
		sharing150_r <= 0;
		sharing151_r <= 0;
		sharing152_r <= 0;
		sharing153_r <= 0;
		sharing154_r <= 0;
		sharing155_r <= 0;
		sharing156_r <= 0;
		sharing157_r <= 0;
		sharing158_r <= 0;
		sharing159_r <= 0;
		sharing160_r <= 0;
		sharing161_r <= 0;
		sharing162_r <= 0;
		sharing163_r <= 0;
		sharing164_r <= 0;
		sharing165_r <= 0;
		sharing166_r <= 0;
		sharing167_r <= 0;
		sharing168_r <= 0;
	end
	else begin
		sharing0_r <= sharing0_w;
		sharing1_r <= sharing1_w;
		sharing2_r <= sharing2_w;
		sharing3_r <= sharing3_w;
		sharing4_r <= sharing4_w;
		sharing5_r <= sharing5_w;
		sharing6_r <= sharing6_w;
		sharing7_r <= sharing7_w;
		sharing8_r <= sharing8_w;
		sharing9_r <= sharing9_w;
		sharing10_r <= sharing10_w;
		sharing11_r <= sharing11_w;
		sharing12_r <= sharing12_w;
		sharing13_r <= sharing13_w;
		sharing14_r <= sharing14_w;
		sharing15_r <= sharing15_w;
		sharing16_r <= sharing16_w;
		sharing17_r <= sharing17_w;
		sharing18_r <= sharing18_w;
		sharing19_r <= sharing19_w;
		sharing20_r <= sharing20_w;
		sharing21_r <= sharing21_w;
		sharing22_r <= sharing22_w;
		sharing23_r <= sharing23_w;
		sharing24_r <= sharing24_w;
		sharing25_r <= sharing25_w;
		sharing26_r <= sharing26_w;
		sharing27_r <= sharing27_w;
		sharing28_r <= sharing28_w;
		sharing29_r <= sharing29_w;
		sharing30_r <= sharing30_w;
		sharing31_r <= sharing31_w;
		sharing32_r <= sharing32_w;
		sharing33_r <= sharing33_w;
		sharing34_r <= sharing34_w;
		sharing35_r <= sharing35_w;
		sharing36_r <= sharing36_w;
		sharing37_r <= sharing37_w;
		sharing38_r <= sharing38_w;
		sharing39_r <= sharing39_w;
		sharing40_r <= sharing40_w;
		sharing41_r <= sharing41_w;
		sharing42_r <= sharing42_w;
		sharing43_r <= sharing43_w;
		sharing44_r <= sharing44_w;
		sharing45_r <= sharing45_w;
		sharing46_r <= sharing46_w;
		sharing47_r <= sharing47_w;
		sharing48_r <= sharing48_w;
		sharing49_r <= sharing49_w;
		sharing50_r <= sharing50_w;
		sharing51_r <= sharing51_w;
		sharing52_r <= sharing52_w;
		sharing53_r <= sharing53_w;
		sharing54_r <= sharing54_w;
		sharing55_r <= sharing55_w;
		sharing56_r <= sharing56_w;
		sharing57_r <= sharing57_w;
		sharing58_r <= sharing58_w;
		sharing59_r <= sharing59_w;
		sharing60_r <= sharing60_w;
		sharing61_r <= sharing61_w;
		sharing62_r <= sharing62_w;
		sharing63_r <= sharing63_w;
		sharing64_r <= sharing64_w;
		sharing65_r <= sharing65_w;
		sharing66_r <= sharing66_w;
		sharing67_r <= sharing67_w;
		sharing68_r <= sharing68_w;
		sharing69_r <= sharing69_w;
		sharing70_r <= sharing70_w;
		sharing71_r <= sharing71_w;
		sharing72_r <= sharing72_w;
		sharing73_r <= sharing73_w;
		sharing74_r <= sharing74_w;
		sharing75_r <= sharing75_w;
		sharing76_r <= sharing76_w;
		sharing77_r <= sharing77_w;
		sharing78_r <= sharing78_w;
		sharing79_r <= sharing79_w;
		sharing80_r <= sharing80_w;
		sharing81_r <= sharing81_w;
		sharing82_r <= sharing82_w;
		sharing83_r <= sharing83_w;
		sharing84_r <= sharing84_w;
		sharing85_r <= sharing85_w;
		sharing86_r <= sharing86_w;
		sharing87_r <= sharing87_w;
		sharing88_r <= sharing88_w;
		sharing89_r <= sharing89_w;
		sharing90_r <= sharing90_w;
		sharing91_r <= sharing91_w;
		sharing92_r <= sharing92_w;
		sharing93_r <= sharing93_w;
		sharing94_r <= sharing94_w;
		sharing95_r <= sharing95_w;
		sharing96_r <= sharing96_w;
		sharing97_r <= sharing97_w;
		sharing98_r <= sharing98_w;
		sharing99_r <= sharing99_w;
		sharing100_r <= sharing100_w;
		sharing101_r <= sharing101_w;
		sharing102_r <= sharing102_w;
		sharing103_r <= sharing103_w;
		sharing104_r <= sharing104_w;
		sharing105_r <= sharing105_w;
		sharing106_r <= sharing106_w;
		sharing107_r <= sharing107_w;
		sharing108_r <= sharing108_w;
		sharing109_r <= sharing109_w;
		sharing110_r <= sharing110_w;
		sharing111_r <= sharing111_w;
		sharing112_r <= sharing112_w;
		sharing113_r <= sharing113_w;
		sharing114_r <= sharing114_w;
		sharing115_r <= sharing115_w;
		sharing116_r <= sharing116_w;
		sharing117_r <= sharing117_w;
		sharing118_r <= sharing118_w;
		sharing119_r <= sharing119_w;
		sharing120_r <= sharing120_w;
		sharing121_r <= sharing121_w;
		sharing122_r <= sharing122_w;
		sharing123_r <= sharing123_w;
		sharing124_r <= sharing124_w;
		sharing125_r <= sharing125_w;
		sharing126_r <= sharing126_w;
		sharing127_r <= sharing127_w;
		sharing128_r <= sharing128_w;
		sharing129_r <= sharing129_w;
		sharing130_r <= sharing130_w;
		sharing131_r <= sharing131_w;
		sharing132_r <= sharing132_w;
		sharing133_r <= sharing133_w;
		sharing134_r <= sharing134_w;
		sharing135_r <= sharing135_w;
		sharing136_r <= sharing136_w;
		sharing137_r <= sharing137_w;
		sharing138_r <= sharing138_w;
		sharing139_r <= sharing139_w;
		sharing140_r <= sharing140_w;
		sharing141_r <= sharing141_w;
		sharing142_r <= sharing142_w;
		sharing143_r <= sharing143_w;
		sharing144_r <= sharing144_w;
		sharing145_r <= sharing145_w;
		sharing146_r <= sharing146_w;
		sharing147_r <= sharing147_w;
		sharing148_r <= sharing148_w;
		sharing149_r <= sharing149_w;
		sharing150_r <= sharing150_w;
		sharing151_r <= sharing151_w;
		sharing152_r <= sharing152_w;
		sharing153_r <= sharing153_w;
		sharing154_r <= sharing154_w;
		sharing155_r <= sharing155_w;
		sharing156_r <= sharing156_w;
		sharing157_r <= sharing157_w;
		sharing158_r <= sharing158_w;
		sharing159_r <= sharing159_w;
		sharing160_r <= sharing160_w;
		sharing161_r <= sharing161_w;
		sharing162_r <= sharing162_w;
		sharing163_r <= sharing163_w;
		sharing164_r <= sharing164_w;
		sharing165_r <= sharing165_w;
		sharing166_r <= sharing166_w;
		sharing167_r <= sharing167_w;
		sharing168_r <= sharing168_w;
	end
end
endmodule
