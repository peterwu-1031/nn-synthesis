module fc1 (
	input [2027:0] in,
	output [127:0] out
);

wire [3:0] relu_out [0:31];
wire [9:0] weighted_sum [0:31];
wire [9:0] sharing0;
wire [9:0] sharing1;
wire [9:0] sharing2;
wire [9:0] sharing3;
wire [9:0] sharing4;
wire [9:0] sharing5;
wire [9:0] sharing6;
wire [9:0] sharing7;
wire [9:0] sharing8;
wire [9:0] sharing9;
wire [9:0] sharing10;
wire [9:0] sharing11;
wire [9:0] sharing12;
wire [9:0] sharing13;
wire [9:0] sharing14;
wire [9:0] sharing15;
wire [9:0] sharing16;
wire [9:0] sharing17;
wire [9:0] sharing18;
wire [9:0] sharing19;
wire [9:0] sharing20;
wire [9:0] sharing21;
wire [9:0] sharing22;
wire [9:0] sharing23;
wire [9:0] sharing24;
wire [9:0] sharing25;
wire [9:0] sharing26;
wire [9:0] sharing27;
wire [9:0] sharing28;
wire [9:0] sharing29;
wire [9:0] sharing30;
wire [9:0] sharing31;
wire [9:0] sharing32;
wire [9:0] sharing33;
wire [9:0] sharing34;
wire [9:0] sharing35;
wire [9:0] sharing36;
wire [9:0] sharing37;
wire [9:0] sharing38;
wire [9:0] sharing39;
wire [9:0] sharing40;
wire [9:0] sharing41;
wire [9:0] sharing42;
wire [9:0] sharing43;
wire [9:0] sharing44;
wire [9:0] sharing45;
wire [9:0] sharing46;
wire [9:0] sharing47;
wire [9:0] sharing48;
wire [9:0] sharing49;
wire [9:0] sharing50;
wire [9:0] sharing51;
wire [9:0] sharing52;
wire [9:0] sharing53;
wire [9:0] sharing54;
wire [9:0] sharing55;
wire [9:0] sharing56;
wire [9:0] sharing57;
wire [9:0] sharing58;
wire [9:0] sharing59;
wire [9:0] sharing60;
wire [9:0] sharing61;
wire [9:0] sharing62;
wire [9:0] sharing63;
wire [9:0] sharing64;
wire [9:0] sharing65;
wire [9:0] sharing66;
wire [9:0] sharing67;
wire [9:0] sharing68;
wire [9:0] sharing69;
wire [9:0] sharing70;
wire [9:0] sharing71;
wire [9:0] sharing72;
wire [9:0] sharing73;
wire [9:0] sharing74;
wire [9:0] sharing75;
wire [9:0] sharing76;
wire [9:0] sharing77;
wire [9:0] sharing78;
wire [9:0] sharing79;
wire [9:0] sharing80;
wire [9:0] sharing81;
wire [9:0] sharing82;
wire [9:0] sharing83;
wire [9:0] sharing84;
wire [9:0] sharing85;
wire [9:0] sharing86;
wire [9:0] sharing87;
wire [9:0] sharing88;
wire [9:0] sharing89;
wire [9:0] sharing90;
wire [9:0] sharing91;
wire [9:0] sharing92;
wire [9:0] sharing93;
wire [9:0] sharing94;
wire [9:0] sharing95;
wire [9:0] sharing96;
wire [9:0] sharing97;
wire [9:0] sharing98;
wire [9:0] sharing99;
wire [9:0] sharing100;
wire [9:0] sharing101;
wire [9:0] sharing102;
wire [9:0] sharing103;
wire [9:0] sharing104;
wire [9:0] sharing105;
wire [9:0] sharing106;
wire [9:0] sharing107;
wire [9:0] sharing108;
wire [9:0] sharing109;
wire [9:0] sharing110;
wire [9:0] sharing111;
wire [9:0] sharing112;
wire [9:0] sharing113;
wire [9:0] sharing114;
wire [9:0] sharing115;
wire [9:0] sharing116;
wire [9:0] sharing117;
wire [9:0] sharing118;
wire [9:0] sharing119;
wire [9:0] sharing120;
wire [9:0] sharing121;
wire [9:0] sharing122;
wire [9:0] sharing123;
wire [9:0] sharing124;
wire [9:0] sharing125;
wire [9:0] sharing126;
wire [9:0] sharing127;
wire [9:0] sharing128;
wire [9:0] sharing129;
wire [9:0] sharing130;
wire [9:0] sharing131;
wire [9:0] sharing132;
wire [9:0] sharing133;
wire [9:0] sharing134;
wire [9:0] sharing135;
wire [9:0] sharing136;
wire [9:0] sharing137;
wire [9:0] sharing138;
wire [9:0] sharing139;
wire [9:0] sharing140;
wire [9:0] sharing141;
wire [9:0] sharing142;
wire [9:0] sharing143;
wire [9:0] sharing144;
wire [9:0] sharing145;
wire [9:0] sharing146;
wire [9:0] sharing147;
wire [9:0] sharing148;
wire [9:0] sharing149;
wire [9:0] sharing150;
wire [9:0] sharing151;
wire [9:0] sharing152;
wire [9:0] sharing153;
wire [9:0] sharing154;
wire [9:0] sharing155;
wire [9:0] sharing156;
wire [9:0] sharing157;
wire [9:0] sharing158;
wire [9:0] sharing159;
wire [9:0] sharing160;
wire [9:0] sharing161;
wire [9:0] sharing162;
wire [9:0] sharing163;
wire [9:0] sharing164;
wire [9:0] sharing165;
wire [9:0] sharing166;
wire [9:0] sharing167;
wire [9:0] sharing168;
wire [9:0] sharing169;
wire [9:0] sharing170;
wire [9:0] sharing171;
wire [9:0] sharing172;
wire [9:0] sharing173;
wire [9:0] sharing174;
wire [9:0] sharing175;
wire [9:0] sharing176;
wire [9:0] sharing177;
wire [9:0] sharing178;
wire [9:0] sharing179;
wire [9:0] sharing180;
wire [9:0] sharing181;
wire [9:0] sharing182;
wire [9:0] sharing183;
wire [9:0] sharing184;
wire [9:0] sharing185;
wire [9:0] sharing186;
wire [9:0] sharing187;
wire [9:0] sharing188;
wire [9:0] sharing189;
wire [9:0] sharing190;
wire [9:0] sharing191;
wire [9:0] sharing192;
wire [9:0] sharing193;
wire [9:0] sharing194;
wire [9:0] sharing195;
wire [9:0] sharing196;
wire [9:0] sharing197;
wire [9:0] sharing198;
wire [9:0] sharing199;
wire [9:0] sharing200;
wire [9:0] sharing201;
wire [9:0] sharing202;
wire [9:0] sharing203;
wire [9:0] sharing204;
wire [9:0] sharing205;
wire [9:0] sharing206;
wire [9:0] sharing207;
wire [9:0] sharing208;
wire [9:0] sharing209;
wire [9:0] sharing210;
wire [9:0] sharing211;
wire [9:0] sharing212;
wire [9:0] sharing213;
wire [9:0] sharing214;
wire [9:0] sharing215;
wire [9:0] sharing216;
wire [9:0] sharing217;
wire [9:0] sharing218;
wire [9:0] sharing219;
wire [9:0] sharing220;
wire [9:0] sharing221;
wire [9:0] sharing222;
wire [9:0] sharing223;
wire [9:0] sharing224;
wire [9:0] sharing225;
wire [9:0] sharing226;
wire [9:0] sharing227;
wire [9:0] sharing228;
wire [9:0] sharing229;
wire [9:0] sharing230;
wire [9:0] sharing231;
wire [9:0] sharing232;
wire [9:0] sharing233;
wire [9:0] sharing234;
wire [9:0] sharing235;
wire [9:0] sharing236;
wire [9:0] sharing237;
wire [9:0] sharing238;
wire [9:0] sharing239;
wire [9:0] sharing240;
wire [9:0] sharing241;
wire [9:0] sharing242;
wire [9:0] sharing243;
wire [9:0] sharing244;
wire [9:0] sharing245;
wire [9:0] sharing246;
wire [9:0] sharing247;
wire [9:0] sharing248;
wire [9:0] sharing249;
wire [9:0] sharing250;
wire [9:0] sharing251;
wire [9:0] sharing252;
wire [9:0] sharing253;
wire [9:0] sharing254;
wire [9:0] sharing255;

assign sharing0 = $signed(in[515-:4])+$signed(in[259-:4])+$signed(in[1795-:4])+$signed(in[1027-:4])+$signed(in[1671-:4])+$signed(in[1287-:4])+$signed(in[1799-:4])+$signed(in[1163-:4])+$signed(in[1291-:4])+$signed(in[655-:4])+$signed(in[271-:4])+$signed(in[1295-:4])+$signed(in[1275-:4])+$signed({in[667-:4],1'b0})+$signed(in[1819-:4])+$signed(in[283-:4])+$signed(in[155-:4])+$signed(in[667-:4])+$signed(in[287-:4])+$signed(in[671-:4])+$signed(in[1279-:4])+$signed(in[935-:4])+$signed({in[1715-:4],1'b0})+$signed(in[1335-:4])+$signed({in[1723-:4],1'b0})+$signed({in[1339-:4],1'b0})+$signed({in[1343-:4],1'b0})+$signed(in[831-:4])+$signed(in[1347-:4])+$signed(in[71-:4])+$signed({in[1611-:4],1'b0})+$signed(in[75-:4])+$signed(in[1739-:4])+$signed(in[331-:4])+$signed({in[975-:4],1'b0})+$signed(in[335-:4])+$signed(in[595-:4])+$signed(in[855-:4])+$signed(in[2007-:4])+$signed(in[1627-:4])+$signed(in[603-:4])+$signed({in[2015-:4],1'b0})+$signed(in[1507-:4])+$signed(in[2019-:4])+$signed({in[615-:4],1'b0})+$signed(in[2023-:4])+$signed(in[875-:4])+$signed(in[379-:4])+$signed(in[247-:4])+$signed(in[251-:4])+$signed({in[1663-:4],1'b0})+$signed(in[1535-:4])+$signed(-in[1415-:4])+$signed(-in[1039-:4])+$signed(-in[527-:4])+$signed(-{in[1427-:4],1'b0})+$signed(-in[795-:4])+$signed(-in[411-:4])+$signed(-in[543-:4])+$signed(-in[799-:4])+$signed(-in[1055-:4])+$signed(-in[547-:4])+$signed(-in[163-:4])+$signed(-in[39-:4])+$signed(-in[1071-:4])+$signed(-in[63-:4])+$signed(-in[1087-:4])+$signed(-in[1091-:4])+$signed(-{in[71-:4],2'b0})+$signed(-in[967-:4])+$signed(-{in[75-:4],2'b0})+$signed(-{in[79-:4],2'b0})+$signed(-in[847-:4])+$signed(-in[1871-:4])+$signed(-{in[95-:4],1'b0})+$signed(-in[363-:4])+$signed(-in[1899-:4])+$signed(-in[751-:4])+$signed(-in[495-:4])+$signed(-in[1139-:4])+$signed(-in[499-:4])+$signed(-in[1019-:4])+$signed(-in[763-:4]);
assign sharing1 = $signed(in[143-:4])+$signed(in[531-:4])+$signed(in[1171-:4])+$signed(in[1175-:4])+$signed(in[1435-:4])+$signed(in[1827-:4])+$signed(in[423-:4])+$signed(in[1831-:4])+$signed(in[427-:4])+$signed({in[1971-:4],1'b0})+$signed(in[1851-:4])+$signed(in[1603-:4])+$signed(in[1879-:4])+$signed(in[1883-:4])+$signed(in[1247-:4])+$signed(in[483-:4])+$signed(in[1763-:4])+$signed(in[1383-:4])+$signed(in[1767-:4])+$signed(in[619-:4])+$signed(in[1259-:4])+$signed(in[2027-:4])+$signed(in[1915-:4])+$signed(-in[519-:4])+$signed(-in[263-:4])+$signed(-in[903-:4])+$signed(-in[1563-:4])+$signed(-in[415-:4])+$signed(-in[1823-:4])+$signed(-in[1311-:4])+$signed(-in[1571-:4])+$signed(-in[167-:4])+$signed(-in[1703-:4])+$signed(-in[179-:4])+$signed(-in[1719-:4])+$signed(-in[955-:4])+$signed(-in[67-:4])+$signed(-in[1107-:4])+$signed(-in[1751-:4])+$signed(-in[91-:4])+$signed(-in[219-:4])+$signed(-in[1755-:4])+$signed(-in[227-:4])+$signed(-in[355-:4])+$signed(-in[111-:4])+$signed(-in[1527-:4]);
assign sharing2 = $signed({in[515-:4],1'b0})+$signed(in[259-:4])+$signed(in[515-:4])+$signed(in[255-:4])+$signed(in[1927-:4])+$signed(in[519-:4])+$signed({in[1931-:4],1'b0})+$signed(in[1803-:4])+$signed(in[1419-:4])+$signed(in[143-:4])+$signed(in[1935-:4])+$signed({in[531-:4],1'b0})+$signed({in[1427-:4],1'b0})+$signed({in[535-:4],1'b0})+$signed(in[1943-:4])+$signed({in[1431-:4],1'b0})+$signed({in[1819-:4],1'b0})+$signed(in[1435-:4])+$signed(in[415-:4])+$signed(in[1951-:4])+$signed({in[1191-:4],1'b0})+$signed(in[1963-:4])+$signed(in[1711-:4])+$signed(in[1715-:4])+$signed(in[307-:4])+$signed(in[1331-:4])+$signed({in[311-:4],1'b0})+$signed(in[1919-:4])+$signed(in[1599-:4])+$signed({in[1475-:4],1'b0})+$signed({in[1479-:4],1'b0})+$signed(in[71-:4])+$signed(in[967-:4])+$signed({in[75-:4],1'b0})+$signed({in[1867-:4],1'b0})+$signed({in[1483-:4],1'b0})+$signed({in[79-:4],1'b0})+$signed(in[79-:4])+$signed(in[207-:4])+$signed(in[1231-:4])+$signed(in[1871-:4])+$signed(in[83-:4])+$signed({in[1487-:4],1'b0})+$signed({in[463-:4],1'b0})+$signed({in[467-:4],1'b0})+$signed(in[1751-:4])+$signed(in[1879-:4])+$signed({in[1491-:4],1'b0})+$signed({in[1243-:4],1'b0})+$signed({in[1883-:4],1'b0})+$signed({in[1495-:4],1'b0})+$signed(in[2007-:4])+$signed(in[987-:4])+$signed(in[1887-:4])+$signed(in[1499-:4])+$signed(in[611-:4])+$signed(in[1763-:4])+$signed(in[1891-:4])+$signed(in[483-:4])+$signed(in[1383-:4])+$signed(in[487-:4])+$signed(in[363-:4])+$signed(in[1899-:4])+$signed(in[1651-:4])+$signed(in[1655-:4])+$signed({in[1915-:4],1'b0})+$signed(in[1531-:4])+$signed({in[511-:4],1'b0})+$signed(in[895-:4])+$signed(-in[1027-:4])+$signed(-in[399-:4])+$signed(-in[407-:4])+$signed(-in[1175-:4])+$signed(-in[1051-:4])+$signed(-in[411-:4])+$signed(-in[1563-:4])+$signed(-in[667-:4])+$signed(-in[1567-:4])+$signed(-in[163-:4])+$signed(-in[167-:4])+$signed(-in[295-:4])+$signed(-in[315-:4])+$signed(-in[319-:4])+$signed(-in[1731-:4])+$signed(-in[1615-:4])+$signed(-in[1103-:4])+$signed(-in[211-:4])+$signed(-in[343-:4])+$signed(-in[1115-:4])+$signed(-in[347-:4])+$signed(-in[351-:4])+$signed(-in[111-:4])+$signed(-in[1775-:4])+$signed(-{in[371-:4],1'b0})+$signed(-in[1271-:4])+$signed(-{in[635-:4],1'b0})+$signed(-in[1787-:4])+$signed(-in[383-:4]);
assign sharing3 = $signed(in[1035-:4])+$signed(in[1107-:4])+$signed(in[1511-:4])+$signed(-in[1347-:4])+$signed(-in[1559-:4])+$signed(-in[455-:4])+$signed(-in[1607-:4])+$signed(-in[2023-:4])+$signed(-in[431-:4])+$signed(-in[1647-:4])+$signed(-in[435-:4])+$signed(-in[819-:4])+$signed(-in[1299-:4])+$signed(-in[1555-:4])+$signed(-in[759-:4])+$signed(-in[1983-:4])+$signed(-in[671-:4]);
assign sharing4 = $signed(in[1027-:4])+$signed(in[1799-:4])+$signed(in[775-:4])+$signed(in[903-:4])+$signed(in[1547-:4])+$signed(in[1803-:4])+$signed(in[399-:4])+$signed(in[1167-:4])+$signed(in[1935-:4])+$signed(in[147-:4])+$signed(in[919-:4])+$signed(in[279-:4])+$signed(in[667-:4])+$signed(in[1695-:4])+$signed(in[671-:4])+$signed(in[799-:4])+$signed(in[1791-:4])+$signed(in[823-:4])+$signed(in[311-:4])+$signed(in[1079-:4])+$signed(in[827-:4])+$signed(in[955-:4])+$signed(in[1731-:4])+$signed(in[327-:4])+$signed({in[1747-:4],1'b0})+$signed(in[851-:4])+$signed(in[859-:4])+$signed(in[91-:4])+$signed(in[1755-:4])+$signed(in[1119-:4])+$signed(in[1503-:4])+$signed(in[871-:4])+$signed(in[1131-:4])+$signed(in[1647-:4])+$signed(in[1651-:4])+$signed(in[1271-:4])+$signed(in[1787-:4])+$signed(in[1663-:4])+$signed(-in[1379-:4])+$signed(-in[1763-:4])+$signed(-in[1767-:4])+$signed(-in[1895-:4])+$signed(-in[71-:4])+$signed(-in[235-:4])+$signed(-in[1967-:4])+$signed(-in[1427-:4])+$signed(-in[1431-:4])+$signed(-in[27-:4])+$signed(-in[31-:4]);
assign sharing5 = $signed(in[899-:4])+$signed(in[1671-:4])+$signed(in[1035-:4])+$signed(in[1679-:4])+$signed(in[527-:4])+$signed(in[275-:4])+$signed(in[539-:4])+$signed(in[1819-:4])+$signed(in[1691-:4])+$signed(in[1439-:4])+$signed(in[163-:4])+$signed(in[931-:4])+$signed(in[1571-:4])+$signed(in[171-:4])+$signed(in[175-:4])+$signed({in[307-:4],1'b0})+$signed(in[1331-:4])+$signed(in[319-:4])+$signed(in[1599-:4])+$signed(in[1855-:4])+$signed(in[1219-:4])+$signed(in[1487-:4])+$signed(in[1871-:4])+$signed({in[1619-:4],1'b0})+$signed(in[467-:4])+$signed(in[979-:4])+$signed(in[2003-:4])+$signed(in[215-:4])+$signed(in[983-:4])+$signed(in[1495-:4])+$signed({in[219-:4],1'b0})+$signed(in[1623-:4])+$signed(in[1627-:4])+$signed(in[1879-:4])+$signed(in[2007-:4])+$signed(in[227-:4])+$signed(in[1891-:4])+$signed(in[487-:4])+$signed(in[1383-:4])+$signed(in[123-:4])+$signed(in[111-:4])+$signed({in[243-:4],1'b0})+$signed(in[1523-:4])+$signed({in[247-:4],1'b0})+$signed({in[1655-:4],1'b0})+$signed({in[1659-:4],1'b0})+$signed(in[251-:4])+$signed({in[255-:4],1'b0})+$signed(in[1535-:4])+$signed(-in[99-:4])+$signed(-in[1059-:4])+$signed(-in[1795-:4])+$signed(-in[1155-:4])+$signed(-in[1123-:4])+$signed(-in[615-:4])+$signed(-in[2027-:4])+$signed(-in[431-:4])+$signed(-in[751-:4])+$signed(-in[1075-:4])+$signed(-in[339-:4])+$signed(-in[1011-:4])+$signed(-in[1139-:4])+$signed(-in[1919-:4])+$signed(-in[767-:4])+$signed(-in[2015-:4])+$signed(-in[763-:4])+$signed(-in[1343-:4]);
assign sharing6 = $signed(in[1667-:4])+$signed(in[659-:4])+$signed(in[663-:4])+$signed({in[667-:4],1'b0})+$signed(in[283-:4])+$signed(in[1691-:4])+$signed({in[1695-:4],1'b0})+$signed(in[163-:4])+$signed(in[291-:4])+$signed(in[803-:4])+$signed(in[1699-:4])+$signed(in[807-:4])+$signed(in[1063-:4])+$signed(in[1191-:4])+$signed(in[1831-:4])+$signed(in[1839-:4])+$signed(in[1663-:4])+$signed(in[1843-:4])+$signed(in[951-:4])+$signed(in[959-:4])+$signed(in[1471-:4])+$signed(in[1599-:4])+$signed(in[1727-:4])+$signed(in[451-:4])+$signed(in[1983-:4])+$signed(in[71-:4])+$signed(in[455-:4])+$signed(in[967-:4])+$signed(in[1607-:4])+$signed(in[75-:4])+$signed(in[463-:4])+$signed(in[1615-:4])+$signed(in[1507-:4])+$signed(in[1767-:4])+$signed(in[1643-:4])+$signed({in[1007-:4],1'b0})+$signed(in[239-:4])+$signed(in[1647-:4])+$signed(in[1775-:4])+$signed(in[1011-:4])+$signed(in[1655-:4])+$signed(in[123-:4])+$signed(in[511-:4])+$signed(-in[615-:4])+$signed(-in[871-:4])+$signed(-in[359-:4])+$signed(-in[1707-:4])+$signed(-in[1963-:4])+$signed(-in[203-:4])+$signed(-in[1295-:4])+$signed(-in[1967-:4])+$signed(-in[591-:4])+$signed(-in[879-:4])+$signed(-in[1971-:4])+$signed(-in[1875-:4])+$signed(-in[883-:4])+$signed(-in[1911-:4])+$signed(-in[1435-:4])+$signed(-in[31-:4])+$signed(-in[543-:4]);
assign sharing7 = $signed(in[1543-:4])+$signed(in[1799-:4])+$signed(in[143-:4])+$signed(in[1935-:4])+$signed(in[275-:4])+$signed(in[1939-:4])+$signed(in[1943-:4])+$signed(in[159-:4])+$signed(in[1567-:4])+$signed(in[1215-:4])+$signed(in[1475-:4])+$signed(in[1479-:4])+$signed(in[1867-:4])+$signed(in[1871-:4])+$signed(in[1623-:4])+$signed(in[215-:4])+$signed(in[1631-:4])+$signed(in[1123-:4])+$signed(in[1635-:4])+$signed(in[1519-:4])+$signed(in[1523-:4])+$signed(-in[771-:4])+$signed(-in[1283-:4])+$signed(-in[775-:4])+$signed(-in[1415-:4])+$signed(-in[1419-:4])+$signed(-in[1423-:4])+$signed(-in[1427-:4])+$signed(-in[27-:4])+$signed(-in[795-:4])+$signed(-in[547-:4])+$signed(-in[1443-:4])+$signed(-in[1827-:4])+$signed(-in[39-:4])+$signed(-in[555-:4])+$signed(-in[827-:4])+$signed(-in[1083-:4])+$signed(-in[63-:4])+$signed(-in[1731-:4])+$signed(-in[335-:4])+$signed(-in[599-:4])+$signed(-in[1879-:4])+$signed(-in[603-:4])+$signed(-in[1883-:4])+$signed(-in[2011-:4])+$signed(-{in[95-:4],1'b0})+$signed(-in[1887-:4])+$signed(-in[867-:4])+$signed(-in[747-:4])+$signed(-in[751-:4])+$signed(-in[1903-:4])+$signed(-in[115-:4])+$signed(-in[759-:4])+$signed(-in[763-:4]);
assign sharing8 = $signed(in[771-:4])+$signed(in[775-:4])+$signed(in[1415-:4])+$signed(in[1803-:4])+$signed(in[403-:4])+$signed(in[1431-:4])+$signed(in[1559-:4])+$signed(in[1531-:4])+$signed({in[411-:4],1'b0})+$signed({in[1819-:4],1'b0})+$signed({in[799-:4],1'b0})+$signed(in[1695-:4])+$signed(in[1951-:4])+$signed(in[1955-:4])+$signed({in[1575-:4],1'b0})+$signed(in[39-:4])+$signed(in[167-:4])+$signed(in[1067-:4])+$signed(in[1079-:4])+$signed(in[1083-:4])+$signed(in[1595-:4])+$signed(in[1087-:4])+$signed(in[1599-:4])+$signed({in[1091-:4],1'b0})+$signed(in[1475-:4])+$signed(in[1479-:4])+$signed({in[75-:4],1'b0})+$signed(in[1483-:4])+$signed(in[1611-:4])+$signed(in[79-:4])+$signed(in[463-:4])+$signed(in[1487-:4])+$signed(in[1615-:4])+$signed(in[1491-:4])+$signed(in[1111-:4])+$signed(in[1751-:4])+$signed({in[91-:4],1'b0})+$signed({in[1499-:4],1'b0})+$signed(in[1627-:4])+$signed(in[1755-:4])+$signed({in[95-:4],1'b0})+$signed(in[1759-:4])+$signed(in[99-:4])+$signed(in[1127-:4])+$signed(in[751-:4])+$signed(in[1015-:4])+$signed(in[759-:4])+$signed(in[1275-:4])+$signed(in[767-:4])+$signed(-in[611-:4])+$signed(-in[423-:4])+$signed(-in[1831-:4])+$signed(-in[2023-:4])+$signed(-in[1927-:4])+$signed(-in[619-:4])+$signed(-in[1211-:4])+$signed(-in[1679-:4])+$signed(-in[1295-:4])+$signed(-in[1967-:4])+$signed(-in[1299-:4])+$signed(-in[563-:4])+$signed(-in[1971-:4])+$signed(-{in[663-:4],1'b0})+$signed(-{in[1687-:4],1'b0})+$signed(-in[1339-:4])+$signed(-in[1723-:4])+$signed(-in[671-:4]);
assign sharing9 = $signed({in[647-:4],1'b0})+$signed(in[519-:4])+$signed(in[651-:4])+$signed(in[1551-:4])+$signed(in[531-:4])+$signed(in[1939-:4])+$signed(in[23-:4])+$signed(in[31-:4])+$signed(in[1311-:4])+$signed(in[1187-:4])+$signed(in[1315-:4])+$signed(in[1319-:4])+$signed(in[1447-:4])+$signed(in[1451-:4])+$signed(in[175-:4])+$signed(in[1327-:4])+$signed(in[947-:4])+$signed(in[1975-:4])+$signed(in[955-:4])+$signed(in[1219-:4])+$signed(in[1603-:4])+$signed(in[199-:4])+$signed(in[1991-:4])+$signed(in[587-:4])+$signed(in[479-:4])+$signed(in[1631-:4])+$signed(in[483-:4])+$signed(in[1379-:4])+$signed(in[231-:4])+$signed(in[999-:4])+$signed(in[235-:4])+$signed(in[1259-:4])+$signed(in[1647-:4])+$signed(in[1915-:4])+$signed(in[511-:4])+$signed(-in[1155-:4])+$signed(-in[391-:4])+$signed(-in[903-:4])+$signed(-in[267-:4])+$signed(-in[151-:4])+$signed(-in[667-:4])+$signed(-in[1835-:4])+$signed(-in[567-:4])+$signed(-in[827-:4])+$signed(-in[1851-:4])+$signed(-in[447-:4])+$signed(-in[1731-:4])+$signed(-in[1607-:4])+$signed(-in[1735-:4])+$signed(-in[331-:4])+$signed(-in[971-:4])+$signed(-in[1739-:4])+$signed(-in[875-:4])+$signed(-in[883-:4])+$signed(-in[1779-:4])+$signed(-in[375-:4])+$signed(-in[1023-:4]);
assign sharing10 = $signed(in[131-:4])+$signed(in[899-:4])+$signed({in[1799-:4],1'b0})+$signed(in[1159-:4])+$signed(in[1031-:4])+$signed(in[1287-:4])+$signed(in[139-:4])+$signed({in[1807-:4],1'b0})+$signed(in[527-:4])+$signed(in[143-:4])+$signed(in[399-:4])+$signed({in[1811-:4],1'b0})+$signed(in[147-:4])+$signed(in[1427-:4])+$signed(in[1431-:4])+$signed(in[1435-:4])+$signed(in[1575-:4])+$signed(in[1579-:4])+$signed(in[555-:4])+$signed(in[1323-:4])+$signed({in[175-:4],1'b0})+$signed(in[435-:4])+$signed(in[1971-:4])+$signed(in[1079-:4])+$signed(in[567-:4])+$signed(in[951-:4])+$signed(in[1339-:4])+$signed({in[1475-:4],1'b0})+$signed({in[1867-:4],1'b0})+$signed(in[75-:4])+$signed(in[1483-:4])+$signed(in[207-:4])+$signed(in[463-:4])+$signed(in[1487-:4])+$signed({in[851-:4],1'b0})+$signed(in[1107-:4])+$signed(in[1235-:4])+$signed(in[467-:4])+$signed({in[1751-:4],1'b0})+$signed(in[1623-:4])+$signed(in[1239-:4])+$signed(in[119-:4])+$signed({in[1755-:4],1'b0})+$signed(in[1243-:4])+$signed({in[1499-:4],1'b0})+$signed(in[2011-:4])+$signed({in[1759-:4],1'b0})+$signed(in[1631-:4])+$signed(in[863-:4])+$signed(in[1635-:4])+$signed(in[2019-:4])+$signed({in[123-:4],1'b0})+$signed(in[1003-:4])+$signed(in[1143-:4])+$signed({in[1915-:4],1'b0})+$signed(in[1787-:4])+$signed(in[1535-:4])+$signed(-in[259-:4])+$signed(-in[1667-:4])+$signed(-{in[263-:4],1'b0})+$signed(-in[1555-:4])+$signed(-in[1563-:4])+$signed(-in[1311-:4])+$signed(-in[287-:4])+$signed(-in[1063-:4])+$signed(-in[1835-:4])+$signed(-in[427-:4])+$signed(-in[303-:4])+$signed(-in[307-:4])+$signed(-in[1719-:4])+$signed(-in[315-:4])+$signed(-in[67-:4])+$signed(-in[1603-:4])+$signed(-in[1987-:4])+$signed(-in[1607-:4])+$signed(-in[1615-:4])+$signed(-in[211-:4])+$signed(-in[987-:4])+$signed(-in[247-:4])+$signed(-in[1647-:4])+$signed(-in[239-:4])+$signed(-in[1263-:4])+$signed(-in[243-:4])+$signed(-in[1655-:4])+$signed(-in[1659-:4])+$signed(-{in[1663-:4],1'b0})+$signed(-in[255-:4]);
assign sharing11 = $signed(in[1059-:4])+$signed(in[1259-:4])+$signed(in[155-:4])+$signed(in[1211-:4])+$signed(in[219-:4])+$signed(in[1711-:4])+$signed(in[1171-:4])+$signed(in[1843-:4])+$signed(in[1619-:4])+$signed(in[635-:4])+$signed(in[1567-:4])+$signed(-in[1827-:4])+$signed(-in[1699-:4])+$signed(-in[1383-:4])+$signed(-in[1831-:4])+$signed(-in[479-:4])+$signed(-in[1131-:4])+$signed(-in[1879-:4])+$signed(-in[1551-:4])+$signed(-in[655-:4])+$signed(-in[431-:4])+$signed(-in[335-:4])+$signed(-in[1015-:4])+$signed(-in[1115-:4])+$signed(-in[1887-:4]);
assign sharing12 = $signed(in[1155-:4])+$signed(in[1671-:4])+$signed(in[907-:4])+$signed(in[1163-:4])+$signed(in[1939-:4])+$signed(in[1051-:4])+$signed(in[543-:4])+$signed(in[927-:4])+$signed({in[1059-:4],1'b0})+$signed(in[1963-:4])+$signed(in[563-:4])+$signed(in[1075-:4])+$signed(in[951-:4])+$signed(in[567-:4])+$signed(in[1207-:4])+$signed(in[315-:4])+$signed(in[571-:4])+$signed(in[583-:4])+$signed(in[967-:4])+$signed(in[1223-:4])+$signed(in[1739-:4])+$signed(in[975-:4])+$signed(in[1743-:4])+$signed(in[1107-:4])+$signed(in[1119-:4])+$signed(in[999-:4])+$signed(in[1271-:4])+$signed({in[1003-:4],1'b0})+$signed({in[1007-:4],1'b0})+$signed(in[1263-:4])+$signed({in[1011-:4],1'b0})+$signed(in[1267-:4])+$signed(in[1911-:4])+$signed(in[635-:4])+$signed(in[1023-:4])+$signed(-in[1927-:4])+$signed(-in[1803-:4])+$signed(-in[1555-:4])+$signed(-in[1659-:4])+$signed(-in[1823-:4])+$signed(-in[1827-:4])+$signed(-in[423-:4])+$signed(-in[1703-:4])+$signed(-in[1707-:4])+$signed(-in[1843-:4])+$signed(-in[1471-:4])+$signed(-in[1475-:4])+$signed(-{in[1739-:4],2'b0})+$signed(-in[335-:4])+$signed(-{in[1747-:4],1'b0})+$signed(-in[343-:4])+$signed(-in[1755-:4])+$signed(-in[479-:4])+$signed(-in[1759-:4])+$signed(-in[883-:4])+$signed(-in[123-:4]);
assign sharing13 = $signed(in[1035-:4])+$signed(in[1167-:4])+$signed(in[1551-:4])+$signed(in[147-:4])+$signed(in[919-:4])+$signed(in[151-:4])+$signed(in[667-:4])+$signed(in[823-:4])+$signed(in[1083-:4])+$signed(in[1723-:4])+$signed(in[191-:4])+$signed(in[1087-:4])+$signed(in[1727-:4])+$signed(in[1347-:4])+$signed(in[1603-:4])+$signed(in[1735-:4])+$signed(in[2015-:4])+$signed(in[2019-:4])+$signed(in[99-:4])+$signed(in[355-:4])+$signed(in[867-:4])+$signed({in[359-:4],1'b0})+$signed(in[1895-:4])+$signed(in[2023-:4])+$signed(in[875-:4])+$signed(in[879-:4])+$signed({in[1783-:4],1'b0})+$signed(in[379-:4])+$signed(in[767-:4])+$signed(-in[391-:4])+$signed(-in[655-:4])+$signed(-in[271-:4])+$signed(-in[279-:4])+$signed(-in[283-:4])+$signed(-in[1567-:4])+$signed(-in[1579-:4])+$signed(-in[1615-:4])+$signed(-in[1871-:4])+$signed(-in[467-:4])+$signed(-in[1623-:4])+$signed(-{in[1627-:4],1'b0})+$signed(-in[347-:4])+$signed(-in[1499-:4])+$signed(-{in[1631-:4],1'b0})+$signed(-in[1763-:4])+$signed(-{in[1767-:4],1'b0})+$signed(-in[231-:4])+$signed(-in[1643-:4]);
assign sharing14 = $signed(in[655-:4])+$signed(in[1807-:4])+$signed({in[1691-:4],1'b0})+$signed(in[1691-:4])+$signed(in[803-:4])+$signed(in[1059-:4])+$signed({in[1727-:4],1'b0})+$signed(in[1727-:4])+$signed(in[1855-:4])+$signed({in[1731-:4],1'b0})+$signed(in[327-:4])+$signed({in[331-:4],1'b0})+$signed(in[335-:4])+$signed(in[863-:4])+$signed({in[1635-:4],1'b0})+$signed(in[867-:4])+$signed(in[1763-:4])+$signed(in[231-:4])+$signed(in[1639-:4])+$signed(in[235-:4])+$signed(in[239-:4])+$signed(in[1519-:4])+$signed(in[371-:4])+$signed(in[1019-:4])+$signed(-{in[1775-:4],1'b0})+$signed(-in[383-:4]);
assign sharing15 = $signed(in[643-:4])+$signed(in[523-:4])+$signed(in[1427-:4])+$signed(in[1431-:4])+$signed({in[1435-:4],1'b0})+$signed({in[1819-:4],1'b0})+$signed(in[923-:4])+$signed(in[1311-:4])+$signed(in[1823-:4])+$signed(in[1439-:4])+$signed(in[35-:4])+$signed(in[1583-:4])+$signed(in[1971-:4])+$signed(in[567-:4])+$signed(in[1467-:4])+$signed(in[1471-:4])+$signed(in[195-:4])+$signed(in[583-:4])+$signed(in[75-:4])+$signed({in[1871-:4],1'b0})+$signed(in[211-:4])+$signed(in[1623-:4])+$signed(in[1627-:4])+$signed(in[479-:4])+$signed(in[1383-:4])+$signed(in[363-:4])+$signed(in[1259-:4])+$signed(in[123-:4])+$signed(in[1263-:4])+$signed(in[1267-:4])+$signed(in[631-:4])+$signed(in[635-:4])+$signed(in[1919-:4])+$signed(-{in[259-:4],1'b0})+$signed(-in[775-:4])+$signed(-in[1551-:4])+$signed(-{in[1687-:4],2'b0})+$signed(-in[663-:4])+$signed(-in[155-:4])+$signed(-in[1051-:4])+$signed(-in[667-:4])+$signed(-{in[287-:4],2'b0})+$signed(-in[1187-:4])+$signed(-in[1191-:4])+$signed(-in[1447-:4])+$signed(-in[827-:4])+$signed(-in[831-:4])+$signed(-{in[323-:4],2'b0})+$signed(-in[1603-:4])+$signed(-{in[207-:4],1'b0})+$signed(-in[1231-:4])+$signed(-in[1747-:4])+$signed(-in[987-:4])+$signed(-in[1499-:4])+$signed(-{in[1503-:4],1'b0})+$signed(-in[999-:4])+$signed(-in[1003-:4])+$signed(-{in[1011-:4],2'b0})+$signed(-in[755-:4])+$signed(-in[883-:4])+$signed(-in[1651-:4])+$signed(-in[1659-:4])+$signed(-in[511-:4]);
assign sharing16 = $signed(in[1539-:4])+$signed(in[515-:4])+$signed(in[1027-:4])+$signed({in[903-:4],1'b0})+$signed(in[647-:4])+$signed(in[1927-:4])+$signed({in[1035-:4],1'b0})+$signed(in[907-:4])+$signed(in[1035-:4])+$signed(in[1807-:4])+$signed(in[1299-:4])+$signed(in[1811-:4])+$signed({in[663-:4],1'b0})+$signed(in[1311-:4])+$signed(in[1315-:4])+$signed(in[1699-:4])+$signed(in[1703-:4])+$signed(in[303-:4])+$signed(in[1075-:4])+$signed({in[951-:4],1'b0})+$signed(in[439-:4])+$signed(in[1079-:4])+$signed(in[1083-:4])+$signed(in[1339-:4])+$signed(in[1347-:4])+$signed(in[1987-:4])+$signed(in[847-:4])+$signed(in[1615-:4])+$signed(in[979-:4])+$signed(in[1107-:4])+$signed(in[1875-:4])+$signed(in[855-:4])+$signed(in[215-:4])+$signed(in[347-:4])+$signed(in[351-:4])+$signed(in[1119-:4])+$signed({in[355-:4],1'b0})+$signed(in[1763-:4])+$signed(in[359-:4])+$signed(in[1127-:4])+$signed(in[1255-:4])+$signed(in[619-:4])+$signed(in[1771-:4])+$signed(in[2027-:4])+$signed(in[623-:4])+$signed({in[1523-:4],1'b0})+$signed(in[1527-:4])+$signed(in[1535-:4])+$signed(-{in[259-:4],1'b0})+$signed(-in[1379-:4])+$signed(-in[1603-:4])+$signed(-in[1559-:4])+$signed(-in[1831-:4])+$signed(-in[1447-:4])+$signed(-in[1643-:4])+$signed(-{in[819-:4],1'b0})+$signed(-in[19-:4])+$signed(-in[83-:4])+$signed(-in[1975-:4])+$signed(-in[1499-:4]);
assign sharing17 = $signed(in[35-:4])+$signed(in[231-:4])+$signed(in[1895-:4])+$signed(in[935-:4])+$signed(in[811-:4])+$signed(in[235-:4])+$signed(in[1455-:4])+$signed(in[1711-:4])+$signed(in[879-:4])+$signed(in[147-:4])+$signed(in[179-:4])+$signed(in[883-:4])+$signed(in[23-:4])+$signed(in[151-:4])+$signed(in[183-:4])+$signed(in[1595-:4])+$signed(in[255-:4])+$signed(-in[1155-:4])+$signed(-in[1667-:4])+$signed(-in[267-:4])+$signed(-in[1039-:4])+$signed(-in[1679-:4])+$signed(-in[919-:4])+$signed(-in[895-:4])+$signed(-{in[1563-:4],1'b0})+$signed(-in[1819-:4])+$signed(-in[803-:4])+$signed(-in[175-:4])+$signed(-in[431-:4])+$signed(-in[307-:4])+$signed(-in[1715-:4])+$signed(-in[1207-:4])+$signed(-in[1851-:4])+$signed(-in[1727-:4])+$signed(-in[1855-:4])+$signed(-in[319-:4])+$signed(-{in[1479-:4],1'b0})+$signed(-in[327-:4])+$signed(-{in[1483-:4],1'b0})+$signed(-in[1739-:4])+$signed(-in[1103-:4])+$signed(-{in[1619-:4],1'b0})+$signed(-in[211-:4])+$signed(-in[467-:4])+$signed(-in[1111-:4])+$signed(-{in[219-:4],1'b0})+$signed(-in[1627-:4])+$signed(-in[223-:4])+$signed(-in[95-:4])+$signed(-in[1631-:4])+$signed(-in[363-:4])+$signed(-in[1515-:4])+$signed(-{in[119-:4],1'b0})+$signed(-in[379-:4])+$signed(-in[127-:4]);
assign sharing18 = $signed(in[891-:4])+$signed(in[1799-:4])+$signed(in[519-:4])+$signed(in[1927-:4])+$signed(in[523-:4])+$signed(in[1931-:4])+$signed(in[1783-:4])+$signed({in[527-:4],1'b0})+$signed(in[1555-:4])+$signed(in[1311-:4])+$signed(in[675-:4])+$signed(in[167-:4])+$signed(in[1319-:4])+$signed(in[1703-:4])+$signed(in[1831-:4])+$signed(in[1711-:4])+$signed(in[1463-:4])+$signed(in[955-:4])+$signed({in[1983-:4],1'b0})+$signed(in[1215-:4])+$signed(in[831-:4])+$signed(in[579-:4])+$signed(in[1219-:4])+$signed(in[1479-:4])+$signed(in[1991-:4])+$signed({in[207-:4],1'b0})+$signed(in[591-:4])+$signed(in[595-:4])+$signed(in[1875-:4])+$signed({in[1879-:4],1'b0})+$signed(in[1503-:4])+$signed(in[483-:4])+$signed(in[1895-:4])+$signed(in[875-:4])+$signed(in[1259-:4])+$signed(in[1771-:4])+$signed(in[1519-:4])+$signed(in[883-:4])+$signed(in[1015-:4])+$signed(in[1523-:4])+$signed(in[1271-:4])+$signed({in[635-:4],1'b0})+$signed(in[507-:4])+$signed({in[1663-:4],1'b0})+$signed(in[383-:4])+$signed(-in[1667-:4])+$signed(-in[263-:4])+$signed(-in[1419-:4])+$signed(-{in[1171-:4],2'b0})+$signed(-in[663-:4])+$signed(-in[1023-:4])+$signed(-in[415-:4])+$signed(-in[299-:4])+$signed(-in[811-:4])+$signed(-{in[431-:4],1'b0})+$signed(-in[447-:4])+$signed(-in[1087-:4])+$signed(-in[67-:4])+$signed(-in[1859-:4])+$signed(-in[971-:4])+$signed(-in[975-:4])+$signed(-in[1103-:4])+$signed(-in[979-:4])+$signed(-in[95-:4])+$signed(-in[99-:4])+$signed(-in[995-:4])+$signed(-in[2027-:4])+$signed(-in[755-:4])+$signed(-in[1651-:4])+$signed(-in[759-:4])+$signed(-in[1659-:4])+$signed(-in[763-:4]);
assign sharing19 = $signed(in[1431-:4])+$signed(in[1819-:4])+$signed(in[1827-:4])+$signed(in[803-:4])+$signed(in[135-:4])+$signed(in[71-:4])+$signed(in[1115-:4])+$signed({in[1775-:4],1'b0})+$signed(in[1679-:4])+$signed(in[79-:4])+$signed(in[1427-:4])+$signed(in[1683-:4])+$signed(in[1467-:4])+$signed(in[83-:4])+$signed(in[1687-:4])+$signed(in[1107-:4])+$signed(in[1111-:4])+$signed(in[1083-:4])+$signed(-in[827-:4])+$signed(-in[1763-:4])+$signed(-in[391-:4])+$signed(-in[1063-:4])+$signed(-in[1067-:4])+$signed(-in[1759-:4])+$signed(-in[659-:4])+$signed(-in[1619-:4])+$signed(-in[215-:4])+$signed(-in[1627-:4])+$signed(-in[1851-:4])+$signed(-in[375-:4])+$signed(-in[767-:4]);
assign sharing20 = $signed(in[1539-:4])+$signed(in[259-:4])+$signed(in[771-:4])+$signed({in[1543-:4],1'b0})+$signed(in[1415-:4])+$signed({in[1547-:4],2'b0})+$signed(in[139-:4])+$signed(in[1035-:4])+$signed({in[1551-:4],1'b0})+$signed(in[1423-:4])+$signed(in[1559-:4])+$signed(in[1435-:4])+$signed(in[1947-:4])+$signed(in[1055-:4])+$signed(in[1059-:4])+$signed(in[1699-:4])+$signed(in[1447-:4])+$signed(in[1327-:4])+$signed(in[307-:4])+$signed(in[1591-:4])+$signed({in[1595-:4],1'b0})+$signed({in[1599-:4],1'b0})+$signed(in[1603-:4])+$signed(in[1987-:4])+$signed(in[1611-:4])+$signed(in[79-:4])+$signed(in[207-:4])+$signed(in[1487-:4])+$signed({in[1491-:4],1'b0})+$signed(in[983-:4])+$signed(in[91-:4])+$signed(in[1115-:4])+$signed(in[1499-:4])+$signed(in[1883-:4])+$signed(in[863-:4])+$signed(in[99-:4])+$signed(in[1891-:4])+$signed(in[359-:4])+$signed(in[1383-:4])+$signed(in[879-:4])+$signed(in[1903-:4])+$signed(in[1663-:4])+$signed(-in[471-:4])+$signed(-in[419-:4])+$signed(-{in[167-:4],1'b0})+$signed(-in[1471-:4])+$signed(-in[847-:4])+$signed(-in[1875-:4])+$signed(-in[115-:4])+$signed(-in[371-:4])+$signed(-in[895-:4])+$signed(-in[1527-:4])+$signed(-in[1723-:4])+$signed(-in[1823-:4]);
assign sharing21 = $signed(in[1155-:4])+$signed(in[907-:4])+$signed(in[911-:4])+$signed({in[1555-:4],1'b0})+$signed(in[147-:4])+$signed(in[155-:4])+$signed({in[931-:4],1'b0})+$signed(in[803-:4])+$signed(in[1571-:4])+$signed({in[935-:4],1'b0})+$signed(in[807-:4])+$signed(in[1191-:4])+$signed(in[1575-:4])+$signed({in[823-:4],1'b0})+$signed(in[311-:4])+$signed(in[1211-:4])+$signed(in[831-:4])+$signed(in[1607-:4])+$signed(in[859-:4])+$signed(in[247-:4])+$signed(in[1507-:4])+$signed(in[759-:4])+$signed(in[375-:4])+$signed(in[251-:4])+$signed(in[255-:4])+$signed(-in[131-:4])+$signed(-in[643-:4])+$signed(-in[1667-:4])+$signed(-in[1671-:4])+$signed(-in[1675-:4])+$signed(-in[271-:4])+$signed(-{in[919-:4],1'b0})+$signed(-in[663-:4])+$signed(-in[1815-:4])+$signed(-in[415-:4])+$signed(-in[291-:4])+$signed(-in[1315-:4])+$signed(-in[947-:4])+$signed(-in[1075-:4])+$signed(-in[1343-:4])+$signed(-in[1091-:4])+$signed(-{in[999-:4],1'b0})+$signed(-in[619-:4])+$signed(-in[1003-:4])+$signed(-in[2027-:4])+$signed(-{in[239-:4],1'b0})+$signed(-in[623-:4])+$signed(-in[1531-:4])+$signed(-{in[639-:4],1'b0});
assign sharing22 = $signed(in[259-:4])+$signed(in[387-:4])+$signed(in[903-:4])+$signed(in[1927-:4])+$signed(in[1655-:4])+$signed({in[1931-:4],1'b0})+$signed(in[1551-:4])+$signed(in[1935-:4])+$signed(in[531-:4])+$signed(in[1555-:4])+$signed(in[1939-:4])+$signed(in[535-:4])+$signed(in[539-:4])+$signed(in[1695-:4])+$signed(in[1187-:4])+$signed(in[1319-:4])+$signed(in[1323-:4])+$signed(in[1327-:4])+$signed(in[1715-:4])+$signed({in[579-:4],1'b0})+$signed(in[1603-:4])+$signed(in[583-:4])+$signed(in[1995-:4])+$signed(in[207-:4])+$signed(in[339-:4])+$signed(in[1747-:4])+$signed(in[1751-:4])+$signed(in[1883-:4])+$signed(in[1887-:4])+$signed(in[1891-:4])+$signed(in[487-:4])+$signed(in[1015-:4])+$signed(in[1019-:4])+$signed({in[1663-:4],1'b0})+$signed(in[511-:4])+$signed(-{in[519-:4],1'b0})+$signed(-in[1035-:4])+$signed(-in[1039-:4])+$signed(-in[1431-:4])+$signed(-in[411-:4])+$signed(-in[1563-:4])+$signed(-in[415-:4])+$signed(-in[803-:4])+$signed(-in[943-:4])+$signed(-in[1847-:4])+$signed(-in[315-:4])+$signed(-in[443-:4])+$signed(-in[319-:4])+$signed(-in[1727-:4])+$signed(-{in[1219-:4],1'b0})+$signed(-in[323-:4])+$signed(-in[71-:4])+$signed(-{in[1867-:4],2'b0})+$signed(-{in[467-:4],1'b0})+$signed(-in[211-:4])+$signed(-in[355-:4])+$signed(-in[995-:4])+$signed(-in[999-:4])+$signed(-in[1767-:4])+$signed(-in[363-:4])+$signed(-in[755-:4])+$signed(-in[759-:4])+$signed(-{in[1919-:4],1'b0});
assign sharing23 = $signed(in[395-:4])+$signed(in[1171-:4])+$signed(in[1055-:4])+$signed(in[427-:4])+$signed(in[431-:4])+$signed(in[1071-:4])+$signed(in[1467-:4])+$signed(in[1723-:4])+$signed(in[1731-:4])+$signed(in[1735-:4])+$signed(in[1871-:4])+$signed(in[343-:4])+$signed(in[1507-:4])+$signed(in[359-:4])+$signed(in[1259-:4])+$signed(in[111-:4])+$signed(in[1263-:4])+$signed(in[115-:4])+$signed(in[1139-:4])+$signed(in[119-:4])+$signed(-in[515-:4])+$signed(-in[1443-:4])+$signed(-in[1447-:4])+$signed(-in[1703-:4])+$signed(-in[1351-:4])+$signed(-in[663-:4])+$signed(-in[823-:4])+$signed(-in[1631-:4])+$signed(-in[847-:4])+$signed(-in[879-:4])+$signed(-in[983-:4])+$signed(-in[979-:4])+$signed(-in[567-:4])+$signed(-in[1499-:4])+$signed(-in[1119-:4])+$signed(-in[255-:4]);
assign sharing24 = $signed(in[647-:4])+$signed({in[1555-:4],1'b0})+$signed(in[1555-:4])+$signed(in[1687-:4])+$signed(in[1559-:4])+$signed(in[1055-:4])+$signed(in[1535-:4])+$signed({in[1583-:4],1'b0})+$signed(in[1967-:4])+$signed({in[1715-:4],1'b0})+$signed(in[179-:4])+$signed(in[567-:4])+$signed(in[1735-:4])+$signed(in[971-:4])+$signed(in[1103-:4])+$signed(in[1491-:4])+$signed(in[1503-:4])+$signed(in[1635-:4])+$signed(in[1263-:4])+$signed(in[1903-:4])+$signed(in[1531-:4])+$signed(in[639-:4])+$signed(-in[439-:4])+$signed(-in[1347-:4])+$signed(-in[1763-:4])+$signed(-in[999-:4])+$signed(-in[2023-:4])+$signed(-in[1031-:4])+$signed(-{in[1003-:4],2'b0})+$signed(-in[1035-:4])+$signed(-in[1419-:4])+$signed(-{in[1007-:4],1'b0})+$signed(-{in[755-:4],1'b0})+$signed(-in[1111-:4]);
assign sharing25 = $signed(in[775-:4])+$signed(in[1547-:4])+$signed(in[663-:4])+$signed(in[155-:4])+$signed(in[31-:4])+$signed(in[671-:4])+$signed(in[1067-:4])+$signed(in[1071-:4])+$signed(in[1075-:4])+$signed(in[823-:4])+$signed(in[1975-:4])+$signed(in[827-:4])+$signed(in[1339-:4])+$signed(in[1599-:4])+$signed(in[1087-:4])+$signed({in[1603-:4],1'b0})+$signed({in[1607-:4],2'b0})+$signed(in[203-:4])+$signed({in[207-:4],1'b0})+$signed(in[1499-:4])+$signed(in[223-:4])+$signed(in[607-:4])+$signed(in[1759-:4])+$signed(in[2015-:4])+$signed(in[1507-:4])+$signed({in[1639-:4],1'b0})+$signed({in[1659-:4],1'b0})+$signed(in[763-:4])+$signed({in[1663-:4],1'b0})+$signed(in[255-:4])+$signed(-in[899-:4])+$signed(-in[1527-:4])+$signed(-in[519-:4])+$signed(-in[523-:4])+$signed(-{in[1427-:4],1'b0})+$signed(-in[895-:4])+$signed(-{in[1435-:4],1'b0})+$signed(-{in[1567-:4],1'b0})+$signed(-in[163-:4])+$signed(-in[1827-:4])+$signed(-in[1915-:4])+$signed(-in[1191-:4])+$signed(-in[427-:4])+$signed(-in[1451-:4])+$signed(-in[1207-:4])+$signed(-in[1467-:4])+$signed(-{in[1475-:4],1'b0})+$signed(-{in[79-:4],1'b0})+$signed(-in[979-:4])+$signed(-in[1875-:4])+$signed(-{in[215-:4],1'b0})+$signed(-in[87-:4])+$signed(-in[219-:4])+$signed(-in[1255-:4])+$signed(-in[1383-:4])+$signed(-in[1767-:4])+$signed(-in[2027-:4])+$signed(-in[1519-:4])+$signed(-in[1775-:4])+$signed(-{in[371-:4],1'b0})+$signed(-in[115-:4])+$signed(-in[1523-:4])+$signed(-in[1779-:4])+$signed(-{in[375-:4],1'b0})+$signed(-in[119-:4])+$signed(-in[123-:4])+$signed(-in[127-:4]);
assign sharing26 = $signed(in[1155-:4])+$signed(in[1923-:4])+$signed({in[519-:4],1'b0})+$signed(in[1159-:4])+$signed(in[1543-:4])+$signed(in[523-:4])+$signed(in[1547-:4])+$signed(in[527-:4])+$signed(in[1423-:4])+$signed(in[1815-:4])+$signed({in[1435-:4],1'b0})+$signed({in[1819-:4],1'b0})+$signed(in[1439-:4])+$signed(in[1063-:4])+$signed(in[431-:4])+$signed(in[1791-:4])+$signed({in[1207-:4],1'b0})+$signed(in[439-:4])+$signed(in[1211-:4])+$signed(in[1215-:4])+$signed(in[1599-:4])+$signed(in[323-:4])+$signed(in[207-:4])+$signed(in[1871-:4])+$signed({in[467-:4],1'b0})+$signed(in[1491-:4])+$signed(in[1111-:4])+$signed(in[1495-:4])+$signed(in[1115-:4])+$signed(in[1243-:4])+$signed(in[1383-:4])+$signed(in[1639-:4])+$signed(in[1259-:4])+$signed(in[1647-:4])+$signed(in[1783-:4])+$signed(in[507-:4])+$signed(in[127-:4])+$signed(-{in[771-:4],1'b0})+$signed(-in[1667-:4])+$signed(-in[1927-:4])+$signed(-in[267-:4])+$signed(-in[275-:4])+$signed(-in[791-:4])+$signed(-in[27-:4])+$signed(-in[1311-:4])+$signed(-in[287-:4])+$signed(-in[39-:4])+$signed(-in[167-:4])+$signed(-in[815-:4])+$signed(-in[1719-:4])+$signed(-{in[1983-:4],1'b0})+$signed(-in[967-:4])+$signed(-in[1615-:4])+$signed(-in[1619-:4])+$signed(-in[343-:4])+$signed(-in[215-:4])+$signed(-in[219-:4])+$signed(-in[223-:4])+$signed(-in[95-:4])+$signed(-in[99-:4])+$signed(-in[359-:4])+$signed(-in[115-:4])+$signed(-in[755-:4])+$signed(-{in[763-:4],1'b0})+$signed(-in[1019-:4])+$signed(-in[1023-:4]);
assign sharing27 = $signed(in[1283-:4])+$signed(in[1551-:4])+$signed(in[147-:4])+$signed({in[151-:4],1'b0})+$signed({in[663-:4],1'b0})+$signed({in[667-:4],1'b0})+$signed(in[1567-:4])+$signed(in[1959-:4])+$signed(in[1707-:4])+$signed(in[1723-:4])+$signed(in[1727-:4])+$signed(in[831-:4])+$signed({in[1347-:4],1'b0})+$signed(in[1235-:4])+$signed(in[1755-:4])+$signed({in[2015-:4],1'b0})+$signed(in[2019-:4])+$signed({in[2023-:4],1'b0})+$signed(in[615-:4])+$signed(in[999-:4])+$signed(in[619-:4])+$signed(in[623-:4])+$signed({in[1011-:4],1'b0})+$signed(-in[643-:4])+$signed(-in[255-:4])+$signed(-in[1163-:4])+$signed(-in[1675-:4])+$signed(-in[1811-:4])+$signed(-in[799-:4])+$signed(-in[803-:4])+$signed(-in[1323-:4])+$signed(-in[1715-:4])+$signed(-in[447-:4])+$signed(-in[63-:4])+$signed(-in[1991-:4])+$signed(-in[1995-:4])+$signed(-in[335-:4])+$signed(-in[1743-:4])+$signed(-in[1999-:4])+$signed(-in[987-:4])+$signed(-in[1635-:4])+$signed(-in[1763-:4])+$signed(-in[631-:4])+$signed(-in[1659-:4])+$signed(-{in[1663-:4],1'b0})+$signed(-in[639-:4]);
assign sharing28 = $signed(in[259-:4])+$signed(in[1795-:4])+$signed(in[1799-:4])+$signed(in[1803-:4])+$signed(in[395-:4])+$signed(in[1423-:4])+$signed(in[19-:4])+$signed({in[1023-:4],1'b0})+$signed(in[919-:4])+$signed(in[151-:4])+$signed(in[895-:4])+$signed(in[1695-:4])+$signed(in[811-:4])+$signed({in[1071-:4],1'b0})+$signed(in[1071-:4])+$signed({in[823-:4],1'b0})+$signed(in[1847-:4])+$signed(in[1219-:4])+$signed(in[1859-:4])+$signed(in[339-:4])+$signed(in[467-:4])+$signed(in[851-:4])+$signed({in[343-:4],1'b0})+$signed({in[95-:4],1'b0})+$signed(in[95-:4])+$signed(in[1631-:4])+$signed({in[99-:4],1'b0})+$signed({in[1123-:4],1'b0})+$signed(in[1635-:4])+$signed(in[1895-:4])+$signed(in[491-:4])+$signed(in[875-:4])+$signed({in[751-:4],1'b0})+$signed(in[1903-:4])+$signed(in[371-:4])+$signed(in[755-:4])+$signed({in[1019-:4],1'b0})+$signed({in[767-:4],1'b0})+$signed(in[767-:4])+$signed(-in[1091-:4])+$signed(-in[1667-:4])+$signed(-in[1383-:4])+$signed(-in[331-:4])+$signed(-in[303-:4])+$signed(-in[1039-:4])+$signed(-in[943-:4])+$signed(-in[1103-:4])+$signed(-in[1647-:4])+$signed(-in[243-:4])+$signed(-in[251-:4])+$signed(-in[663-:4])+$signed(-in[1563-:4])+$signed(-in[959-:4])+$signed(-in[123-:4])+$signed(-in[1087-:4]);
assign sharing29 = $signed(in[643-:4])+$signed(in[647-:4])+$signed(in[1927-:4])+$signed(in[1655-:4])+$signed(in[267-:4])+$signed(in[139-:4])+$signed(in[651-:4])+$signed(in[1419-:4])+$signed(in[143-:4])+$signed(in[287-:4])+$signed(in[1823-:4])+$signed(in[1567-:4])+$signed(in[419-:4])+$signed(in[1187-:4])+$signed(in[1315-:4])+$signed(in[295-:4])+$signed(in[1191-:4])+$signed(in[1319-:4])+$signed(in[1703-:4])+$signed(in[999-:4])+$signed(in[1143-:4])+$signed(in[635-:4])+$signed(-in[387-:4])+$signed(-in[1299-:4])+$signed(-in[1171-:4])+$signed(-{in[1559-:4],1'b0})+$signed(-in[1815-:4])+$signed(-in[1175-:4])+$signed(-{in[1819-:4],1'b0})+$signed(-{in[1971-:4],1'b0})+$signed(-in[1715-:4])+$signed(-in[1343-:4])+$signed(-in[451-:4])+$signed(-in[1347-:4])+$signed(-in[1351-:4])+$signed(-in[1607-:4])+$signed(-in[1863-:4])+$signed(-in[203-:4])+$signed(-in[1611-:4])+$signed(-in[1739-:4])+$signed(-{in[2023-:4],1'b0})+$signed(-in[1127-:4])+$signed(-in[2027-:4])+$signed(-in[623-:4])+$signed(-in[1659-:4]);
assign sharing30 = $signed(in[1027-:4])+$signed(in[899-:4])+$signed(in[1927-:4])+$signed(in[1031-:4])+$signed(in[531-:4])+$signed({in[1819-:4],1'b0})+$signed(in[1435-:4])+$signed({in[1567-:4],1'b0})+$signed(in[1311-:4])+$signed(in[1823-:4])+$signed(in[1571-:4])+$signed(in[163-:4])+$signed(in[931-:4])+$signed(in[1575-:4])+$signed(in[167-:4])+$signed(in[1831-:4])+$signed(in[1067-:4])+$signed(in[1851-:4])+$signed(in[1467-:4])+$signed(in[451-:4])+$signed(in[1987-:4])+$signed(in[1479-:4])+$signed(in[971-:4])+$signed({in[975-:4],1'b0})+$signed(in[1103-:4])+$signed(in[1743-:4])+$signed(in[1871-:4])+$signed({in[979-:4],1'b0})+$signed(in[1107-:4])+$signed(in[1875-:4])+$signed({in[983-:4],1'b0})+$signed(in[475-:4])+$signed(in[1503-:4])+$signed({in[1515-:4],1'b0})+$signed(in[1771-:4])+$signed(in[1263-:4])+$signed(in[1775-:4])+$signed(in[1519-:4])+$signed(in[499-:4])+$signed({in[247-:4],1'b0})+$signed(in[895-:4])+$signed(-{in[771-:4],1'b0})+$signed(-in[1415-:4])+$signed(-in[1547-:4])+$signed(-in[1419-:4])+$signed(-in[1039-:4])+$signed(-in[911-:4])+$signed(-{in[1555-:4],2'b0})+$signed(-in[19-:4])+$signed(-in[147-:4])+$signed(-in[659-:4])+$signed(-in[1299-:4])+$signed(-in[23-:4])+$signed(-in[279-:4])+$signed(-in[27-:4])+$signed(-in[671-:4])+$signed(-in[803-:4])+$signed(-in[1443-:4])+$signed(-in[39-:4])+$signed(-in[807-:4])+$signed(-in[1447-:4])+$signed(-in[43-:4])+$signed(-in[1195-:4])+$signed(-in[811-:4])+$signed(-in[1451-:4])+$signed(-in[815-:4])+$signed(-in[567-:4])+$signed(-in[823-:4])+$signed(-in[827-:4])+$signed(-in[63-:4])+$signed(-in[831-:4])+$signed(-in[67-:4])+$signed(-in[327-:4])+$signed(-in[75-:4])+$signed(-in[855-:4])+$signed(-in[1495-:4])+$signed(-in[1371-:4])+$signed(-in[1499-:4])+$signed(-{in[1503-:4],2'b0})+$signed(-{in[95-:4],1'b0})+$signed(-in[1247-:4])+$signed(-in[1375-:4])+$signed(-in[747-:4])+$signed(-{in[751-:4],1'b0})+$signed(-{in[755-:4],1'b0})+$signed(-{in[759-:4],1'b0})+$signed(-in[1143-:4])+$signed(-{in[763-:4],1'b0})+$signed(-{in[767-:4],1'b0})+$signed(-in[127-:4]);
assign sharing31 = $signed(in[1539-:4])+$signed(in[1671-:4])+$signed(in[907-:4])+$signed(in[271-:4])+$signed(in[403-:4])+$signed(in[791-:4])+$signed(in[407-:4])+$signed(in[1659-:4])+$signed(in[1055-:4])+$signed(in[1183-:4])+$signed(in[1711-:4])+$signed(in[1839-:4])+$signed(in[1207-:4])+$signed(in[1083-:4])+$signed(in[1723-:4])+$signed(in[319-:4])+$signed(in[1087-:4])+$signed(in[959-:4])+$signed(in[323-:4])+$signed(in[1603-:4])+$signed(in[211-:4])+$signed(in[987-:4])+$signed(in[631-:4])+$signed(in[1131-:4])+$signed(in[1135-:4])+$signed(in[379-:4])+$signed(in[1139-:4])+$signed(in[503-:4])+$signed(in[635-:4])+$signed(-in[1635-:4])+$signed(-in[287-:4])+$signed(-in[391-:4])+$signed(-in[199-:4])+$signed(-in[1639-:4])+$signed(-in[663-:4])+$signed(-in[203-:4])+$signed(-in[1167-:4])+$signed(-in[919-:4])+$signed(-in[1943-:4])+$signed(-in[1171-:4])+$signed(-in[443-:4])+$signed(-in[599-:4])+$signed(-in[1115-:4])+$signed(-in[1691-:4])+$signed(-in[1119-:4]);
assign sharing32 = $signed({in[259-:4],1'b0})+$signed({in[1539-:4],1'b0})+$signed({in[1675-:4],1'b0})+$signed({in[1551-:4],1'b0})+$signed(in[1807-:4])+$signed({in[659-:4],1'b0})+$signed(in[1939-:4])+$signed({in[663-:4],1'b0})+$signed({in[1559-:4],1'b0})+$signed(in[1051-:4])+$signed({in[927-:4],1'b0})+$signed({in[935-:4],1'b0})+$signed(in[295-:4])+$signed(in[299-:4])+$signed(in[943-:4])+$signed({in[1591-:4],1'b0})+$signed(in[1723-:4])+$signed({in[1599-:4],1'b0})+$signed(in[959-:4])+$signed(in[195-:4])+$signed(in[451-:4])+$signed({in[1607-:4],1'b0})+$signed(in[1483-:4])+$signed({in[207-:4],1'b0})+$signed({in[979-:4],1'b0})+$signed(in[479-:4])+$signed({in[1647-:4],1'b0})+$signed(-in[1859-:4])+$signed(-in[523-:4])+$signed(-in[1419-:4])+$signed(-in[1423-:4])+$signed(-{in[755-:4],1'b0})+$signed(-in[1907-:4])+$signed(-in[1911-:4])+$signed(-in[1083-:4])+$signed(-in[343-:4])+$signed(-in[159-:4]);
assign sharing33 = $signed(in[559-:4])+$signed(in[1963-:4])+$signed(in[1211-:4])+$signed(in[1015-:4])+$signed(-in[1463-:4])+$signed(-in[267-:4])+$signed(-in[535-:4])+$signed(-in[1983-:4])+$signed(-{in[1567-:4],1'b0})+$signed(-in[351-:4]);
assign sharing34 = $signed(in[1283-:4])+$signed(in[1539-:4])+$signed(in[135-:4])+$signed(in[1543-:4])+$signed(in[1959-:4])+$signed(in[1547-:4])+$signed(in[1483-:4])+$signed(in[607-:4])+$signed(in[559-:4])+$signed(in[1999-:4])+$signed(in[2003-:4])+$signed(in[883-:4])+$signed(in[599-:4])+$signed(in[1279-:4])+$signed(-in[471-:4])+$signed(-in[1667-:4])+$signed(-in[1223-:4])+$signed(-in[623-:4])+$signed(-{in[1079-:4],1'b0})+$signed(-in[631-:4])+$signed(-{in[1083-:4],1'b0});
assign sharing35 = $signed(in[1863-:4])+$signed(in[303-:4])+$signed(in[1911-:4])+$signed(in[1875-:4])+$signed(in[1527-:4])+$signed(in[1627-:4])+$signed(in[475-:4])+$signed(in[1759-:4])+$signed(-in[919-:4])+$signed(-{in[1067-:4],1'b0})+$signed(-in[971-:4])+$signed(-in[767-:4]);
assign sharing36 = $signed(in[1863-:4])+$signed(in[71-:4])+$signed(in[1931-:4])+$signed({in[527-:4],1'b0})+$signed(in[847-:4])+$signed(in[1879-:4])+$signed(in[1907-:4])+$signed(in[1911-:4])+$signed(in[571-:4])+$signed({in[1631-:4],1'b0})+$signed(in[959-:4])+$signed(-{in[771-:4],1'b0})+$signed(-{in[935-:4],2'b0})+$signed(-in[1415-:4])+$signed(-{in[1611-:4],2'b0})+$signed(-in[307-:4])+$signed(-{in[1559-:4],2'b0})+$signed(-in[23-:4])+$signed(-{in[283-:4],1'b0})+$signed(-in[311-:4])+$signed(-in[1375-:4]);
assign sharing37 = $signed(in[1671-:4])+$signed(in[1675-:4])+$signed(in[1739-:4])+$signed(in[1783-:4])+$signed(-in[2019-:4])+$signed(-in[263-:4])+$signed(-in[623-:4])+$signed(-in[815-:4])+$signed(-in[1011-:4])+$signed(-in[951-:4])+$signed(-in[1119-:4]);
assign sharing38 = $signed(in[1315-:4])+$signed(in[1539-:4])+$signed(in[1643-:4])+$signed(in[1579-:4])+$signed(in[1327-:4])+$signed(in[979-:4])+$signed(in[319-:4])+$signed(-in[291-:4])+$signed(-in[103-:4])+$signed(-in[551-:4])+$signed(-in[895-:4])+$signed(-in[759-:4])+$signed(-in[1375-:4]);
assign sharing39 = $signed({in[643-:4],2'b0})+$signed({in[647-:4],2'b0})+$signed({in[651-:4],2'b0})+$signed({in[655-:4],2'b0})+$signed(in[279-:4])+$signed(in[1711-:4])+$signed({in[1335-:4],1'b0})+$signed({in[1987-:4],1'b0})+$signed(in[1607-:4])+$signed(in[587-:4])+$signed(in[203-:4])+$signed({in[599-:4],1'b0})+$signed({in[2007-:4],1'b0})+$signed({in[607-:4],1'b0})+$signed(in[611-:4])+$signed(in[867-:4])+$signed(in[879-:4])+$signed(in[1007-:4])+$signed(in[883-:4])+$signed(-in[1891-:4])+$signed(-in[675-:4])+$signed(-in[1475-:4])+$signed(-in[1863-:4])+$signed(-in[135-:4])+$signed(-in[487-:4])+$signed(-in[1895-:4])+$signed(-in[1835-:4])+$signed(-in[1195-:4])+$signed(-in[1867-:4])+$signed(-in[1003-:4])+$signed(-in[1855-:4])+$signed(-in[1143-:4])+$signed(-in[1887-:4]);
assign sharing40 = $signed({in[135-:4],1'b0})+$signed(in[1639-:4])+$signed(in[135-:4])+$signed(in[235-:4])+$signed(in[1579-:4])+$signed({in[1583-:4],1'b0})+$signed(in[655-:4])+$signed({in[1587-:4],1'b0})+$signed(in[83-:4])+$signed(in[535-:4])+$signed(in[183-:4])+$signed(in[1627-:4])+$signed(in[1051-:4])+$signed(in[1207-:4])+$signed(-in[199-:4])+$signed(-in[875-:4])+$signed(-in[791-:4]);
assign sharing41 = $signed(in[579-:4])+$signed(in[231-:4])+$signed(in[423-:4])+$signed(in[631-:4])+$signed(in[523-:4])+$signed(in[175-:4])+$signed(in[819-:4])+$signed(in[855-:4])+$signed(-in[1431-:4])+$signed(-{in[531-:4],1'b0})+$signed(-{in[1495-:4],1'b0})+$signed(-in[87-:4])+$signed(-in[1919-:4]);
assign sharing42 = $signed(in[131-:4])+$signed(in[1623-:4])+$signed({in[1867-:4],1'b0})+$signed(in[1003-:4])+$signed(in[1707-:4])+$signed(in[1879-:4])+$signed(in[1263-:4])+$signed(in[1519-:4])+$signed(in[119-:4])+$signed(in[1271-:4])+$signed({in[123-:4],1'b0})+$signed(in[795-:4])+$signed(in[415-:4])+$signed(-in[1287-:4])+$signed(-{in[1611-:4],2'b0})+$signed(-in[1291-:4])+$signed(-in[815-:4])+$signed(-in[311-:4])+$signed(-in[1659-:4])+$signed(-{in[1663-:4],1'b0});
assign sharing43 = $signed(in[1443-:4])+$signed(in[27-:4])+$signed(in[1547-:4])+$signed(in[43-:4])+$signed(in[1387-:4])+$signed(in[543-:4])+$signed(in[1651-:4])+$signed(in[1655-:4])+$signed(in[1371-:4])+$signed(in[1375-:4])+$signed(-{in[323-:4],1'b0})+$signed(-in[1511-:4])+$signed(-in[295-:4])+$signed(-in[1031-:4])+$signed(-{in[271-:4],1'b0})+$signed(-in[1775-:4])+$signed(-{in[979-:4],1'b0})+$signed(-in[1171-:4])+$signed(-{in[983-:4],1'b0})+$signed(-in[1815-:4])+$signed(-in[1051-:4])+$signed(-in[1823-:4]);
assign sharing44 = $signed(in[1215-:4])+$signed({in[1795-:4],1'b0})+$signed(in[1155-:4])+$signed({in[1767-:4],1'b0})+$signed(in[1991-:4])+$signed(in[1163-:4])+$signed(in[1931-:4])+$signed(in[1995-:4])+$signed(in[363-:4])+$signed(in[1999-:4])+$signed(in[1815-:4])+$signed(in[1847-:4])+$signed({in[1471-:4],1'b0})+$signed(in[1023-:4])+$signed(-in[1543-:4])+$signed(-in[231-:4])+$signed(-{in[1651-:4],1'b0})+$signed(-in[1587-:4])+$signed(-in[311-:4])+$signed(-{in[667-:4],1'b0})+$signed(-in[375-:4]);
assign sharing45 = $signed(in[775-:4])+$signed(in[71-:4])+$signed(in[2023-:4])+$signed(in[1707-:4])+$signed(in[1423-:4])+$signed({in[819-:4],1'b0})+$signed(in[83-:4])+$signed(in[151-:4])+$signed(in[859-:4])+$signed(-in[1267-:4])+$signed(-in[1223-:4]);
assign sharing46 = $signed({in[1859-:4],1'b0})+$signed(in[1027-:4])+$signed(in[963-:4])+$signed({in[1863-:4],1'b0})+$signed(in[1687-:4])+$signed(in[1967-:4])+$signed(in[819-:4])+$signed(in[1919-:4])+$signed(in[1111-:4])+$signed(in[407-:4])+$signed({in[959-:4],1'b0})+$signed(in[383-:4])+$signed(-in[339-:4])+$signed(-in[1451-:4])+$signed(-in[63-:4]);
assign sharing47 = $signed(in[811-:4])+$signed(in[623-:4])+$signed(in[495-:4])+$signed(in[671-:4])+$signed(in[1779-:4])+$signed(in[639-:4])+$signed(-in[1883-:4])+$signed(-in[579-:4])+$signed(-in[1439-:4])+$signed(-in[1675-:4])+$signed(-in[171-:4])+$signed(-in[1771-:4])+$signed(-in[1231-:4])+$signed(-in[1583-:4])+$signed(-in[503-:4])+$signed(-in[1819-:4])+$signed(-in[1335-:4])+$signed(-in[1183-:4]);
assign sharing48 = $signed(in[1571-:4])+$signed(in[963-:4])+$signed({in[487-:4],1'b0})+$signed(in[1351-:4])+$signed(in[171-:4])+$signed(in[587-:4])+$signed(in[1167-:4])+$signed(in[111-:4])+$signed(in[1275-:4])+$signed(in[1983-:4])+$signed(-{in[1767-:4],1'b0})+$signed(-{in[1159-:4],1'b0})+$signed(-in[75-:4])+$signed(-{in[1871-:4],1'b0})+$signed(-in[1423-:4])+$signed(-in[1435-:4])+$signed(-in[799-:4])+$signed(-{in[1211-:4],1'b0})+$signed(-in[315-:4])+$signed(-in[1919-:4]);
assign sharing49 = $signed(in[1867-:4])+$signed({in[1031-:4],1'b0})+$signed(-{in[1507-:4],1'b0})+$signed(-in[1795-:4])+$signed(-in[583-:4])+$signed(-{in[1611-:4],1'b0})+$signed(-in[1195-:4])+$signed(-in[1847-:4])+$signed(-in[1011-:4])+$signed(-in[1143-:4])+$signed(-in[1755-:4]);
assign sharing50 = $signed({in[1827-:4],1'b0})+$signed(in[1743-:4])+$signed({in[1207-:4],1'b0})+$signed(in[183-:4])+$signed({in[475-:4],1'b0})+$signed(in[155-:4])+$signed(in[1691-:4])+$signed({in[1823-:4],1'b0})+$signed(in[639-:4])+$signed(-{in[1059-:4],1'b0})+$signed(-in[771-:4])+$signed(-{in[1091-:4],1'b0})+$signed(-in[1623-:4])+$signed(-in[1575-:4])+$signed(-{in[1107-:4],2'b0})+$signed(-in[247-:4])+$signed(-in[571-:4])+$signed(-{in[379-:4],1'b0})+$signed(-in[923-:4]);
assign sharing51 = $signed(in[1159-:4])+$signed(in[1163-:4])+$signed({in[1167-:4],1'b0})+$signed({in[311-:4],1'b0})+$signed(in[667-:4])+$signed(in[1791-:4])+$signed(-{in[1115-:4],1'b0})+$signed(-in[1643-:4])+$signed(-in[1699-:4])+$signed(-in[463-:4]);
assign sharing52 = $signed(in[99-:4])+$signed(in[1795-:4])+$signed(in[295-:4])+$signed(in[1803-:4])+$signed(in[1551-:4])+$signed(in[1791-:4])+$signed(in[1983-:4])+$signed(in[923-:4])+$signed(in[1663-:4])+$signed(-{in[71-:4],1'b0})+$signed(-in[779-:4])+$signed(-{in[1423-:4],1'b0})+$signed(-in[851-:4])+$signed(-in[915-:4]);
assign sharing53 = $signed({in[259-:4],1'b0})+$signed(in[1379-:4])+$signed(in[615-:4])+$signed({in[1611-:4],1'b0})+$signed(in[1679-:4])+$signed(in[1295-:4])+$signed(in[1683-:4])+$signed(in[563-:4])+$signed({in[311-:4],1'b0})+$signed(in[1655-:4])+$signed(in[1243-:4])+$signed(in[863-:4])+$signed(-{in[1667-:4],1'b0})+$signed(-{in[263-:4],1'b0})+$signed(-{in[267-:4],1'b0})+$signed(-in[1807-:4])+$signed(-in[1811-:4])+$signed(-{in[1815-:4],1'b0})+$signed(-{in[1563-:4],1'b0})+$signed(-in[1179-:4])+$signed(-in[415-:4])+$signed(-in[159-:4])+$signed(-in[431-:4])+$signed(-in[1719-:4])+$signed(-in[955-:4])+$signed(-in[315-:4])+$signed(-in[1855-:4])+$signed(-in[1859-:4])+$signed(-in[455-:4])+$signed(-in[1511-:4])+$signed(-in[1015-:4])+$signed(-in[507-:4]);
assign sharing54 = $signed(in[439-:4])+$signed(in[867-:4])+$signed(in[1635-:4])+$signed(in[387-:4])+$signed(in[963-:4])+$signed(in[455-:4])+$signed(in[855-:4])+$signed(in[755-:4])+$signed(in[87-:4])+$signed(in[791-:4])+$signed(in[383-:4])+$signed(-{in[1635-:4],2'b0})+$signed(-in[579-:4])+$signed(-{in[583-:4],1'b0})+$signed(-in[1931-:4])+$signed(-{in[1263-:4],1'b0})+$signed(-{in[1715-:4],1'b0})+$signed(-in[179-:4])+$signed(-in[183-:4])+$signed(-in[127-:4]);
assign sharing55 = $signed(in[359-:4])+$signed(in[935-:4])+$signed(in[1867-:4])+$signed(in[1567-:4])+$signed(in[495-:4])+$signed(in[1039-:4])+$signed(in[927-:4])+$signed(-in[67-:4])+$signed(-in[1347-:4])+$signed(-in[1579-:4])+$signed(-in[623-:4])+$signed(-in[915-:4]);
assign sharing56 = $signed(in[827-:4])+$signed(in[515-:4])+$signed(in[487-:4])+$signed(in[871-:4])+$signed(in[71-:4])+$signed(in[39-:4])+$signed(in[43-:4])+$signed(in[1451-:4])+$signed(in[75-:4])+$signed(in[747-:4])+$signed(in[1899-:4])+$signed({in[819-:4],1'b0})+$signed({in[755-:4],1'b0})+$signed(in[1759-:4])+$signed({in[91-:4],1'b0})+$signed(in[1243-:4])+$signed(in[1119-:4])+$signed(-in[263-:4])+$signed(-in[2015-:4]);
assign sharing57 = $signed({in[579-:4],1'b0})+$signed(in[583-:4])+$signed(in[967-:4])+$signed({in[971-:4],1'b0})+$signed(in[1291-:4])+$signed(in[843-:4])+$signed(in[1515-:4])+$signed(in[1007-:4])+$signed(in[1523-:4])+$signed({in[1983-:4],1'b0})+$signed(in[1023-:4])+$signed(-{in[1603-:4],1'b0})+$signed(-{in[1663-:4],1'b0})+$signed(-in[1163-:4])+$signed(-{in[307-:4],1'b0})+$signed(-in[275-:4])+$signed(-in[1555-:4])+$signed(-in[1107-:4])+$signed(-in[1975-:4])+$signed(-{in[987-:4],1'b0})+$signed(-{in[255-:4],1'b0})+$signed(-in[351-:4]);
assign sharing58 = $signed({in[1187-:4],1'b0})+$signed(in[67-:4])+$signed({in[1183-:4],1'b0})+$signed({in[1835-:4],1'b0})+$signed(in[651-:4])+$signed(in[1195-:4])+$signed({in[459-:4],1'b0})+$signed(in[1371-:4])+$signed(in[1143-:4])+$signed(in[503-:4])+$signed(in[1659-:4])+$signed({in[479-:4],1'b0})+$signed(in[1535-:4])+$signed(-in[323-:4])+$signed(-in[227-:4])+$signed(-in[395-:4])+$signed(-in[271-:4])+$signed(-in[1619-:4])+$signed(-in[1111-:4])+$signed(-in[1079-:4])+$signed(-in[219-:4])+$signed(-in[279-:4]);
assign sharing59 = $signed(in[195-:4])+$signed({in[1163-:4],1'b0})+$signed(in[587-:4])+$signed(in[1167-:4])+$signed(in[847-:4])+$signed(in[439-:4])+$signed(in[443-:4])+$signed(in[1439-:4])+$signed(-in[963-:4])+$signed(-in[427-:4])+$signed(-in[1135-:4])+$signed(-in[403-:4])+$signed(-in[1463-:4])+$signed(-in[1339-:4])+$signed(-in[1087-:4])+$signed(-in[1055-:4]);
assign sharing60 = $signed(in[1159-:4])+$signed(in[1867-:4])+$signed({in[1743-:4],1'b0})+$signed(in[1807-:4])+$signed(in[815-:4])+$signed(in[759-:4])+$signed(in[1791-:4])+$signed(-in[291-:4])+$signed(-in[35-:4])+$signed(-in[1463-:4])+$signed(-in[1015-:4]);
assign sharing61 = $signed(in[1891-:4])+$signed({in[391-:4],2'b0})+$signed({in[1799-:4],1'b0})+$signed(in[439-:4])+$signed(in[799-:4])+$signed(-in[159-:4])+$signed(-in[163-:4])+$signed(-in[1987-:4])+$signed(-in[995-:4])+$signed(-{in[263-:4],1'b0})+$signed(-in[1719-:4])+$signed(-in[239-:4])+$signed(-in[367-:4])+$signed(-in[531-:4])+$signed(-in[211-:4])+$signed(-in[1619-:4])+$signed(-in[631-:4])+$signed(-{in[1311-:4],1'b0})+$signed(-in[255-:4]);
assign sharing62 = $signed(in[515-:4])+$signed({in[1003-:4],1'b0})+$signed(in[331-:4])+$signed({in[1643-:4],1'b0})+$signed(in[1843-:4])+$signed({in[319-:4],1'b0})+$signed(in[1055-:4])+$signed(-in[1571-:4])+$signed(-in[1987-:4])+$signed(-in[1319-:4])+$signed(-in[471-:4])+$signed(-in[91-:4]);
assign sharing63 = $signed({in[1683-:4],1'b0})+$signed(in[811-:4])+$signed(in[411-:4])+$signed(in[1687-:4])+$signed(-in[1347-:4])+$signed(-in[871-:4])+$signed(-in[2023-:4])+$signed(-in[427-:4])+$signed(-in[911-:4])+$signed(-in[283-:4])+$signed(-in[1975-:4])+$signed(-{in[571-:4],1'b0})+$signed(-in[379-:4])+$signed(-in[191-:4]);
assign sharing64 = $signed(in[1343-:4])+$signed({in[2023-:4],1'b0})+$signed(in[1735-:4])+$signed(in[1611-:4])+$signed({in[1167-:4],1'b0})+$signed({in[1487-:4],1'b0})+$signed(in[983-:4])+$signed(in[115-:4])+$signed(in[243-:4])+$signed(in[1971-:4])+$signed(in[663-:4])+$signed(in[923-:4])+$signed(in[375-:4])+$signed(-in[1135-:4])+$signed(-in[915-:4])+$signed(-{in[759-:4],1'b0})+$signed(-{in[767-:4],1'b0})+$signed(-in[1407-:4]);
assign sharing65 = $signed(in[563-:4])+$signed(in[827-:4])+$signed(in[79-:4])+$signed(-{in[899-:4],1'b0})+$signed(-{in[1575-:4],1'b0})+$signed(-in[999-:4])+$signed(-{in[171-:4],1'b0})+$signed(-{in[1467-:4],1'b0})+$signed(-in[1531-:4]);
assign sharing66 = $signed(in[1603-:4])+$signed(in[99-:4])+$signed(in[1955-:4])+$signed(in[915-:4])+$signed(in[1019-:4])+$signed(-in[1219-:4]);
assign sharing67 = $signed(in[391-:4])+$signed(in[1159-:4])+$signed(in[139-:4])+$signed(in[1487-:4])+$signed(in[1071-:4])+$signed(in[251-:4])+$signed(in[539-:4])+$signed(in[1755-:4])+$signed(-{in[1059-:4],1'b0})+$signed(-in[1127-:4])+$signed(-{in[1131-:4],1'b0})+$signed(-in[1179-:4])+$signed(-{in[1135-:4],1'b0})+$signed(-{in[1783-:4],1'b0})+$signed(-in[23-:4])+$signed(-in[379-:4]);
assign sharing68 = $signed(in[1607-:4])+$signed({in[275-:4],1'b0})+$signed({in[959-:4],1'b0})+$signed(in[279-:4])+$signed(-in[619-:4])+$signed(-in[819-:4]);
assign sharing69 = $signed({in[579-:4],1'b0})+$signed({in[423-:4],1'b0})+$signed({in[1927-:4],1'b0})+$signed({in[83-:4],1'b0})+$signed(in[1815-:4])+$signed(in[1979-:4])+$signed({in[1983-:4],1'b0})+$signed(-{in[99-:4],1'b0})+$signed(-{in[1671-:4],2'b0})+$signed(-in[759-:4])+$signed(-in[1711-:4])+$signed(-in[1335-:4])+$signed(-{in[95-:4],1'b0})+$signed(-in[799-:4]);
assign sharing70 = $signed(in[1739-:4])+$signed(in[1839-:4])+$signed(in[435-:4])+$signed(in[1847-:4])+$signed(in[1471-:4])+$signed(-in[547-:4])+$signed(-in[1603-:4])+$signed(-in[1511-:4])+$signed(-in[1291-:4])+$signed(-{in[271-:4],1'b0})+$signed(-in[155-:4]);
assign sharing71 = $signed(in[875-:4])+$signed(in[635-:4])+$signed(in[1751-:4])+$signed(-in[1883-:4])+$signed(-in[131-:4])+$signed(-{in[1479-:4],1'b0})+$signed(-in[1191-:4])+$signed(-in[75-:4])+$signed(-in[563-:4])+$signed(-in[603-:4])+$signed(-{in[1631-:4],1'b0});
assign sharing72 = $signed({in[643-:4],1'b0})+$signed({in[647-:4],1'b0})+$signed(in[1575-:4])+$signed(in[371-:4])+$signed({in[375-:4],1'b0})+$signed(in[1335-:4])+$signed(in[891-:4])+$signed(in[639-:4])+$signed(-{in[67-:4],1'b0})+$signed(-in[619-:4])+$signed(-in[1163-:4])+$signed(-in[2023-:4]);
assign sharing73 = $signed(in[287-:4])+$signed(-in[483-:4])+$signed(-{in[847-:4],1'b0})+$signed(-{in[851-:4],1'b0})+$signed(-in[595-:4])+$signed(-in[1243-:4])+$signed(-in[415-:4]);
assign sharing74 = $signed(in[803-:4])+$signed(in[1763-:4])+$signed(in[227-:4])+$signed({in[359-:4],1'b0})+$signed(in[1191-:4])+$signed(in[807-:4])+$signed(in[1643-:4])+$signed({in[79-:4],1'b0})+$signed({in[83-:4],1'b0})+$signed({in[1523-:4],1'b0})+$signed({in[1495-:4],1'b0})+$signed({in[1527-:4],1'b0})+$signed(in[1179-:4])+$signed({in[127-:4],1'b0})+$signed(in[1471-:4])+$signed(-in[1727-:4])+$signed(-in[379-:4])+$signed(-in[1715-:4])+$signed(-in[975-:4]);
assign sharing75 = $signed(in[583-:4])+$signed(-{in[1163-:4],1'b0})+$signed(-in[1795-:4])+$signed(-in[559-:4]);
assign sharing76 = $signed({in[803-:4],1'b0})+$signed(in[771-:4])+$signed(in[1123-:4])+$signed(in[615-:4])+$signed(in[871-:4])+$signed(in[523-:4])+$signed(in[491-:4])+$signed(in[1291-:4])+$signed(in[751-:4])+$signed(in[1907-:4])+$signed(in[1947-:4])+$signed(in[1855-:4])+$signed(-{in[659-:4],1'b0})+$signed(-in[1559-:4])+$signed(-{in[1695-:4],1'b0})+$signed(-in[1983-:4]);
assign sharing77 = $signed(in[1283-:4])+$signed(in[1731-:4])+$signed(in[607-:4])+$signed(in[603-:4])+$signed(in[127-:4])+$signed(-in[1091-:4])+$signed(-in[327-:4])+$signed(-in[23-:4])+$signed(-{in[1723-:4],1'b0})+$signed(-in[187-:4])+$signed(-{in[319-:4],1'b0});
assign sharing78 = $signed(in[1859-:4])+$signed(in[227-:4])+$signed(in[519-:4])+$signed(in[431-:4])+$signed(in[1523-:4])+$signed(in[1531-:4])+$signed(in[1211-:4])+$signed(-{in[1711-:4],1'b0})+$signed(-in[1695-:4]);
assign sharing79 = $signed(in[1379-:4])+$signed(in[935-:4])+$signed(in[1511-:4])+$signed(in[1611-:4])+$signed(in[83-:4])+$signed(in[947-:4])+$signed(in[375-:4])+$signed(in[1887-:4])+$signed(-in[1683-:4])+$signed(-in[1063-:4])+$signed(-in[95-:4]);
assign sharing80 = $signed({in[1611-:4],1'b0})+$signed({in[207-:4],1'b0})+$signed(in[495-:4])+$signed({in[883-:4],1'b0})+$signed(in[567-:4])+$signed({in[1499-:4],1'b0})+$signed(in[763-:4])+$signed({in[1503-:4],1'b0})+$signed(-in[1479-:4])+$signed(-in[1519-:4])+$signed(-in[1615-:4])+$signed(-in[315-:4])+$signed(-in[319-:4]);
assign sharing81 = $signed(in[299-:4])+$signed(in[1427-:4])+$signed(in[335-:4])+$signed(in[1439-:4])+$signed(-in[1123-:4])+$signed(-in[1923-:4])+$signed(-in[1767-:4])+$signed(-in[1931-:4])+$signed(-in[571-:4]);
assign sharing82 = $signed(in[407-:4])+$signed({in[1987-:4],1'b0})+$signed({in[643-:4],1'b0})+$signed(in[419-:4])+$signed({in[1315-:4],1'b0})+$signed(in[1511-:4])+$signed(in[1003-:4])+$signed(in[791-:4])+$signed(in[951-:4])+$signed(in[947-:4])+$signed(in[1559-:4])+$signed({in[1787-:4],1'b0})+$signed({in[671-:4],1'b0})+$signed(in[479-:4])+$signed(-in[1923-:4])+$signed(-{in[427-:4],2'b0})+$signed(-in[619-:4])+$signed(-in[1967-:4])+$signed(-in[1495-:4]);
assign sharing83 = $signed(in[1815-:4])+$signed(in[287-:4])+$signed(-in[1299-:4]);
assign sharing84 = $signed(in[291-:4])+$signed(in[1219-:4])+$signed(in[1799-:4])+$signed(in[1211-:4])+$signed(in[879-:4])+$signed(in[339-:4])+$signed(in[1747-:4])+$signed(in[1019-:4])+$signed(-in[1455-:4])+$signed(-in[1407-:4]);
assign sharing85 = $signed(in[227-:4])+$signed(in[1699-:4])+$signed(in[1703-:4])+$signed(in[1611-:4])+$signed(in[1003-:4])+$signed({in[1559-:4],1'b0})+$signed(in[1751-:4])+$signed(in[1787-:4])+$signed(-in[423-:4])+$signed(-in[1159-:4])+$signed(-in[843-:4])+$signed(-{in[847-:4],1'b0})+$signed(-in[975-:4]);
assign sharing86 = $signed(in[1859-:4])+$signed(in[1115-:4])+$signed(-{in[571-:4],1'b0})+$signed(-in[1691-:4])+$signed(-{in[311-:4],1'b0})+$signed(-in[1215-:4]);
assign sharing87 = $signed(in[931-:4])+$signed({in[807-:4],1'b0})+$signed(in[71-:4])+$signed(in[139-:4])+$signed({in[815-:4],1'b0})+$signed(in[207-:4])+$signed({in[851-:4],1'b0})+$signed({in[823-:4],1'b0})+$signed({in[1815-:4],1'b0})+$signed(in[763-:4])+$signed({in[415-:4],1'b0})+$signed(in[1503-:4])+$signed(-{in[1547-:4],1'b0})+$signed(-in[1663-:4])+$signed(-{in[1543-:4],1'b0})+$signed(-in[639-:4]);
assign sharing88 = $signed(in[1239-:4])+$signed(in[1955-:4])+$signed(in[1287-:4])+$signed(in[511-:4])+$signed(-in[931-:4])+$signed(-in[403-:4])+$signed(-{in[311-:4],1'b0});
assign sharing89 = $signed({in[67-:4],1'b0})+$signed({in[291-:4],1'b0})+$signed(in[1415-:4])+$signed(in[1575-:4])+$signed(in[1747-:4])+$signed({in[759-:4],1'b0})+$signed(in[23-:4])+$signed(in[1499-:4])+$signed(in[1467-:4])+$signed(in[1691-:4])+$signed(-in[1431-:4])+$signed(-{in[1871-:4],1'b0})+$signed(-in[1295-:4])+$signed(-in[1591-:4])+$signed(-in[1535-:4]);
assign sharing90 = $signed(in[871-:4])+$signed(in[1287-:4])+$signed(in[203-:4])+$signed({in[147-:4],1'b0})+$signed({in[563-:4],1'b0})+$signed(in[1235-:4])+$signed({in[1939-:4],1'b0})+$signed({in[1239-:4],1'b0})+$signed({in[91-:4],1'b0})+$signed(in[1979-:4])+$signed({in[1947-:4],1'b0})+$signed(in[127-:4])+$signed(-in[1155-:4])+$signed(-in[1031-:4])+$signed(-{in[263-:4],1'b0})+$signed(-in[1023-:4]);
assign sharing91 = $signed({in[811-:4],1'b0})+$signed(in[1903-:4])+$signed(in[1423-:4])+$signed(in[1907-:4])+$signed({in[1975-:4],1'b0})+$signed(in[1211-:4])+$signed({in[1215-:4],1'b0});
assign sharing92 = $signed(in[659-:4])+$signed(in[1631-:4])+$signed(-in[463-:4])+$signed(-in[407-:4])+$signed(-in[1239-:4])+$signed(-in[475-:4])+$signed(-in[511-:4]);
assign sharing93 = $signed({in[1923-:4],1'b0})+$signed(in[35-:4])+$signed(in[767-:4])+$signed(in[23-:4])+$signed(in[31-:4])+$signed(-in[1159-:4])+$signed(-in[171-:4])+$signed(-in[1967-:4])+$signed(-in[1103-:4])+$signed(-in[2003-:4])+$signed(-in[119-:4])+$signed(-in[927-:4]);
assign sharing94 = $signed({in[423-:4],1'b0})+$signed(in[1127-:4])+$signed(in[1607-:4])+$signed(in[1835-:4])+$signed(in[847-:4])+$signed(in[399-:4])+$signed(in[371-:4])+$signed({in[1883-:4],1'b0})+$signed(in[1531-:4])+$signed({in[479-:4],1'b0})+$signed(-{in[1707-:4],1'b0})+$signed(-{in[1711-:4],2'b0})+$signed(-in[1071-:4]);
assign sharing95 = $signed(in[943-:4])+$signed(in[411-:4])+$signed({in[303-:4],1'b0})+$signed(in[1175-:4])+$signed(-in[539-:4])+$signed(-in[543-:4]);
assign sharing96 = $signed({in[611-:4],1'b0})+$signed({in[1543-:4],2'b0})+$signed({in[1547-:4],1'b0})+$signed({in[1491-:4],1'b0})+$signed(in[1695-:4])+$signed(-in[43-:4])+$signed(-in[27-:4]);
assign sharing97 = $signed(in[1651-:4])+$signed(in[1691-:4])+$signed({in[311-:4],1'b0})+$signed(in[1975-:4])+$signed(-in[1035-:4])+$signed(-in[1875-:4])+$signed(-in[347-:4])+$signed(-in[1479-:4]);
assign sharing98 = $signed({in[1571-:4],1'b0})+$signed(in[1315-:4])+$signed(in[931-:4])+$signed({in[1575-:4],1'b0})+$signed(-in[831-:4])+$signed(-in[1343-:4]);
assign sharing99 = $signed({in[75-:4],1'b0})+$signed({in[1479-:4],1'b0})+$signed(in[1423-:4])+$signed(-{in[963-:4],1'b0})+$signed(-in[235-:4]);
assign sharing100 = $signed(in[839-:4])+$signed(in[1515-:4])+$signed(in[651-:4])+$signed(in[427-:4])+$signed(in[1995-:4])+$signed(in[879-:4])+$signed(in[1999-:4])+$signed({in[155-:4],1'b0})+$signed(-in[1091-:4])+$signed(-in[363-:4])+$signed(-in[1863-:4]);
assign sharing101 = $signed(in[1887-:4])+$signed(in[807-:4])+$signed(-in[515-:4]);
assign sharing102 = $signed(in[1319-:4])+$signed(in[1111-:4])+$signed(in[583-:4]);
assign sharing103 = $signed(in[1727-:4])+$signed(in[1667-:4])+$signed({in[663-:4],2'b0})+$signed(in[207-:4]);
assign sharing104 = $signed({in[131-:4],1'b0})+$signed(in[263-:4])+$signed(in[459-:4])+$signed(in[1595-:4])+$signed(in[1723-:4])+$signed({in[127-:4],1'b0})+$signed(-in[1447-:4])+$signed(-in[567-:4]);
assign sharing105 = $signed(in[1987-:4])+$signed(in[1835-:4])+$signed(in[1003-:4])+$signed(in[1779-:4])+$signed(in[1139-:4])+$signed(-in[563-:4])+$signed(-in[899-:4])+$signed(-in[551-:4]);
assign sharing106 = $signed(in[1467-:4])+$signed(in[1543-:4])+$signed(in[1987-:4])+$signed(in[1063-:4]);
assign sharing107 = $signed(in[1667-:4])+$signed(in[1947-:4])+$signed({in[1639-:4],1'b0})+$signed(in[1195-:4])+$signed({in[1583-:4],1'b0})+$signed({in[535-:4],1'b0})+$signed(in[1563-:4])+$signed(-in[2019-:4])+$signed(-in[907-:4])+$signed(-in[335-:4])+$signed(-in[1843-:4])+$signed(-in[987-:4])+$signed(-in[831-:4]);
assign sharing108 = $signed(in[1859-:4])+$signed(in[391-:4])+$signed(in[123-:4])+$signed(in[1683-:4])+$signed(in[1627-:4])+$signed(in[571-:4])+$signed(-in[1139-:4])+$signed(-in[1823-:4]);
assign sharing109 = $signed(in[1463-:4])+$signed(in[903-:4])+$signed({in[1071-:4],1'b0})+$signed(in[855-:4])+$signed(in[1343-:4])+$signed(-in[647-:4])+$signed(-in[483-:4])+$signed(-in[651-:4])+$signed(-in[1671-:4]);
assign sharing110 = $signed({in[1923-:4],1'b0})+$signed({in[1867-:4],1'b0})+$signed(in[2027-:4])+$signed(in[559-:4])+$signed(in[1107-:4])+$signed({in[375-:4],1'b0})+$signed(in[955-:4])+$signed(in[1247-:4])+$signed(-{in[1703-:4],1'b0})+$signed(-in[303-:4])+$signed(-{in[339-:4],1'b0})+$signed(-{in[1655-:4],1'b0})+$signed(-in[1183-:4]);
assign sharing111 = $signed(in[795-:4])+$signed(in[899-:4])+$signed(-in[1779-:4]);
assign sharing112 = $signed(in[1827-:4])+$signed({in[143-:4],1'b0})+$signed({in[83-:4],1'b0})+$signed(in[179-:4])+$signed(in[467-:4])+$signed({in[87-:4],1'b0})+$signed(-in[1719-:4])+$signed(-{in[267-:4],1'b0})+$signed(-in[367-:4])+$signed(-{in[215-:4],1'b0})+$signed(-in[1783-:4]);
assign sharing113 = $signed(in[1727-:4])+$signed(-in[1247-:4])+$signed(-{in[1263-:4],1'b0})+$signed(-in[287-:4]);
assign sharing114 = $signed(in[579-:4])+$signed(in[1843-:4])+$signed({in[1879-:4],1'b0})+$signed(in[1463-:4])+$signed({in[635-:4],1'b0})+$signed({in[1983-:4],1'b0})+$signed(-in[2015-:4])+$signed(-in[1895-:4])+$signed(-in[799-:4]);
assign sharing115 = $signed(in[335-:4])+$signed(in[1239-:4])+$signed(-in[1063-:4])+$signed(-in[2027-:4])+$signed(-{in[1103-:4],1'b0})+$signed(-{in[1615-:4],1'b0})+$signed(-in[927-:4]);
assign sharing116 = $signed({in[1731-:4],1'b0})+$signed({in[1739-:4],1'b0})+$signed(in[1123-:4])+$signed(in[1695-:4])+$signed(-in[103-:4]);
assign sharing117 = $signed(in[643-:4])+$signed(in[1715-:4])+$signed(-in[467-:4])+$signed(-in[1039-:4])+$signed(-in[475-:4])+$signed(-in[1471-:4]);
assign sharing118 = $signed(in[1223-:4])+$signed(in[1767-:4])+$signed(in[1863-:4])+$signed(in[1159-:4])+$signed(in[1163-:4])+$signed(in[1871-:4])+$signed(in[1463-:4])+$signed(in[1175-:4])+$signed(in[1055-:4])+$signed(-in[1243-:4]);
assign sharing119 = $signed(in[499-:4])+$signed(in[863-:4])+$signed(-{in[659-:4],1'b0})+$signed(-in[1923-:4])+$signed(-{in[1983-:4],1'b0})+$signed(-{in[635-:4],1'b0});
assign sharing120 = $signed(in[1851-:4])+$signed(in[1707-:4])+$signed({in[1015-:4],1'b0})+$signed(in[983-:4])+$signed(in[443-:4])+$signed(in[1755-:4])+$signed(-in[175-:4])+$signed(-in[1587-:4])+$signed(-in[31-:4]);
assign sharing121 = $signed({in[1827-:4],1'b0})+$signed(in[1991-:4])+$signed({in[1931-:4],1'b0})+$signed(in[1771-:4])+$signed({in[1879-:4],1'b0})+$signed(in[215-:4])+$signed(in[27-:4])+$signed(in[63-:4])+$signed(-{in[935-:4],1'b0});
assign sharing122 = $signed(in[91-:4])+$signed(in[1611-:4])+$signed(in[1275-:4])+$signed(-{in[1027-:4],1'b0})+$signed(-in[1763-:4])+$signed(-in[267-:4])+$signed(-{in[1075-:4],1'b0})+$signed(-in[347-:4])+$signed(-in[351-:4]);
assign sharing123 = $signed(in[331-:4])+$signed(in[1899-:4])+$signed({in[1175-:4],1'b0})+$signed(in[499-:4])+$signed(-in[1115-:4])+$signed(-in[931-:4]);
assign sharing124 = $signed({in[1171-:4],1'b0})+$signed(in[1915-:4])+$signed(in[971-:4])+$signed(in[1215-:4])+$signed(-in[463-:4])+$signed(-in[891-:4])+$signed(-in[987-:4])+$signed(-in[2007-:4]);
assign sharing125 = $signed({in[1847-:4],1'b0})+$signed(in[1507-:4])+$signed({in[1791-:4],1'b0})+$signed(-in[1255-:4])+$signed(-in[1323-:4])+$signed(-in[1327-:4]);
assign sharing126 = $signed(in[1587-:4])+$signed({in[667-:4],1'b0})+$signed(in[635-:4])+$signed(in[1071-:4])+$signed(-in[675-:4])+$signed(-{in[871-:4],1'b0})+$signed(-{in[879-:4],2'b0})+$signed(-{in[883-:4],2'b0})+$signed(-{in[827-:4],1'b0})+$signed(-{in[1663-:4],2'b0})+$signed(-{in[1759-:4],1'b0});
assign sharing127 = $signed(in[771-:4])+$signed(in[1635-:4])+$signed(in[1555-:4])+$signed(in[1991-:4])+$signed(-{in[1475-:4],1'b0})+$signed(-{in[1579-:4],1'b0})+$signed(-in[1431-:4]);
assign sharing128 = $signed(in[199-:4])+$signed(in[995-:4])+$signed(in[1063-:4])+$signed(in[1471-:4])+$signed(-in[1583-:4]);
assign sharing129 = $signed(in[1707-:4])+$signed(in[1327-:4])+$signed(in[175-:4])+$signed(in[1587-:4])+$signed(in[147-:4])+$signed(-in[803-:4])+$signed(-in[451-:4])+$signed(-in[1839-:4]);
assign sharing130 = $signed(in[1163-:4])+$signed({in[1871-:4],1'b0})+$signed(in[983-:4])+$signed(-in[1643-:4])+$signed(-in[1691-:4])+$signed(-in[1267-:4]);
assign sharing131 = $signed({in[167-:4],1'b0})+$signed(in[1319-:4])+$signed({in[303-:4],1'b0})+$signed({in[655-:4],1'b0})+$signed(in[1327-:4])+$signed(in[947-:4])+$signed({in[855-:4],1'b0});
assign sharing132 = $signed(in[2015-:4])+$signed(in[1595-:4])+$signed(in[1187-:4])+$signed(in[911-:4]);
assign sharing133 = $signed(in[371-:4])+$signed(in[631-:4])+$signed(-{in[1907-:4],1'b0})+$signed(-in[1747-:4])+$signed(-{in[1903-:4],1'b0})+$signed(-{in[1815-:4],1'b0});
assign sharing134 = $signed({in[1931-:4],1'b0})+$signed(in[551-:4])+$signed(in[1935-:4])+$signed(-in[1027-:4])+$signed(-in[303-:4]);
assign sharing135 = $signed({in[1891-:4],1'b0})+$signed(in[547-:4])+$signed({in[1039-:4],1'b0})+$signed({in[87-:4],1'b0})+$signed(in[1883-:4])+$signed(in[1439-:4])+$signed(-{in[259-:4],1'b0});
assign sharing136 = $signed({in[1195-:4],1'b0})+$signed({in[1963-:4],1'b0})+$signed({in[1967-:4],1'b0})+$signed({in[563-:4],1'b0})+$signed({in[1911-:4],1'b0})+$signed({in[2011-:4],1'b0})+$signed(in[1119-:4])+$signed(-in[419-:4]);
assign sharing137 = $signed({in[1803-:4],1'b0})+$signed(in[395-:4])+$signed(-in[1775-:4])+$signed(-{in[671-:4],1'b0})+$signed(-in[959-:4]);
assign sharing138 = $signed(in[159-:4])+$signed(in[67-:4])+$signed({in[1767-:4],1'b0})+$signed(in[627-:4])+$signed(in[1875-:4])+$signed(in[415-:4])+$signed(-in[1371-:4])+$signed(-in[1339-:4])+$signed(-in[1699-:4])+$signed(-in[751-:4]);
assign sharing139 = $signed(in[1651-:4])+$signed(in[979-:4])+$signed(in[1551-:4])+$signed(-in[527-:4])+$signed(-in[607-:4]);
assign sharing140 = $signed(in[355-:4])+$signed({in[147-:4],1'b0})+$signed(in[1819-:4])+$signed(-{in[1311-:4],1'b0})+$signed(-in[1511-:4]);
assign sharing141 = $signed({in[1611-:4],1'b0})+$signed(in[1831-:4])+$signed(-{in[1667-:4],1'b0})+$signed(-in[1083-:4])+$signed(-in[1523-:4]);
assign sharing142 = $signed(-{in[487-:4],2'b0})+$signed(-{in[1863-:4],1'b0})+$signed(-in[875-:4])+$signed(-in[1295-:4])+$signed(-in[495-:4])+$signed(-{in[1971-:4],1'b0})+$signed(-in[1215-:4]);
assign sharing143 = $signed({in[1103-:4],1'b0})+$signed({in[1063-:4],1'b0})+$signed(in[1407-:4])+$signed(-in[1527-:4]);
assign sharing144 = $signed(in[1571-:4])+$signed(in[1799-:4])+$signed(in[1787-:4])+$signed(in[1495-:4])+$signed(-{in[1247-:4],1'b0})+$signed(-in[1999-:4]);
assign sharing145 = $signed({in[95-:4],1'b0})+$signed(in[143-:4])+$signed(-in[423-:4]);
assign sharing146 = $signed(in[167-:4])+$signed(in[587-:4])+$signed({in[591-:4],1'b0})+$signed({in[595-:4],1'b0})+$signed({in[1943-:4],1'b0})+$signed(in[543-:4])+$signed(-in[403-:4])+$signed(-in[447-:4]);
assign sharing147 = $signed(in[1035-:4])+$signed(in[115-:4])+$signed(in[1211-:4])+$signed(in[87-:4])+$signed(-{in[1035-:4],2'b0})+$signed(-in[279-:4]);
assign sharing148 = $signed(in[1855-:4])+$signed(in[775-:4])+$signed(-in[1547-:4])+$signed(-in[1131-:4]);
assign sharing149 = $signed(in[1859-:4])+$signed({in[967-:4],1'b0})+$signed({in[1451-:4],1'b0})+$signed(in[1067-:4])+$signed({in[287-:4],1'b0})+$signed(in[1375-:4])+$signed(-in[923-:4]);
assign sharing150 = $signed(in[987-:4])+$signed(in[151-:4])+$signed(-in[1379-:4])+$signed(-in[363-:4])+$signed(-in[1263-:4]);
assign sharing151 = $signed({in[235-:4],1'b0})+$signed(in[1075-:4])+$signed({in[915-:4],1'b0})+$signed(-in[1563-:4])+$signed(-in[139-:4]);
assign sharing152 = $signed({in[1507-:4],1'b0})+$signed(in[275-:4])+$signed(in[1647-:4])+$signed(-in[1883-:4]);
assign sharing153 = $signed(in[587-:4])+$signed(in[427-:4])+$signed(in[459-:4])+$signed(in[251-:4]);
assign sharing154 = $signed({in[1787-:4],1'b0})+$signed(in[351-:4])+$signed({in[1775-:4],1'b0})+$signed(in[1079-:4])+$signed(-in[1951-:4]);
assign sharing155 = $signed({in[883-:4],1'b0})+$signed({in[1679-:4],1'b0})+$signed(in[327-:4])+$signed(-{in[1515-:4],1'b0})+$signed(-in[1987-:4]);
assign sharing156 = $signed({in[379-:4],1'b0})+$signed({in[1007-:4],1'b0})+$signed(-in[259-:4])+$signed(-in[263-:4])+$signed(-{in[1711-:4],1'b0})+$signed(-in[971-:4]);
assign sharing157 = $signed(in[747-:4])+$signed(in[1735-:4])+$signed(-in[607-:4]);
assign sharing158 = $signed({in[635-:4],2'b0})+$signed(in[1547-:4])+$signed({in[639-:4],1'b0})+$signed(in[1591-:4])+$signed(-in[611-:4])+$signed(-{in[1959-:4],1'b0})+$signed(-{in[895-:4],1'b0})+$signed(-{in[859-:4],1'b0})+$signed(-{in[863-:4],1'b0});
assign sharing159 = $signed(in[487-:4])+$signed({in[755-:4],1'b0})+$signed(in[1419-:4])+$signed(in[1455-:4])+$signed(-{in[1691-:4],1'b0})+$signed(-in[155-:4])+$signed(-{in[935-:4],1'b0});
assign sharing160 = $signed({in[1635-:4],1'b0})+$signed(in[1699-:4])+$signed(-{in[371-:4],1'b0});
assign sharing161 = $signed(in[1731-:4])+$signed(in[1155-:4])+$signed(in[1791-:4])+$signed(in[1559-:4])+$signed(in[639-:4])+$signed(-in[99-:4]);
assign sharing162 = $signed(in[1891-:4])+$signed(-{in[987-:4],1'b0})+$signed(-{in[1055-:4],1'b0});
assign sharing163 = $signed(-in[1487-:4])+$signed(-in[867-:4])+$signed(-in[631-:4])+$signed(-in[455-:4]);
assign sharing164 = $signed({in[199-:4],1'b0})+$signed({in[1703-:4],1'b0})+$signed({in[1707-:4],1'b0})+$signed({in[875-:4],1'b0})+$signed({in[1651-:4],1'b0})+$signed(in[1491-:4])+$signed({in[151-:4],1'b0})+$signed({in[251-:4],1'b0})+$signed(-in[411-:4])+$signed(-in[1111-:4]);
assign sharing165 = $signed(in[291-:4])+$signed(in[763-:4])+$signed({in[375-:4],1'b0})+$signed(in[1311-:4])+$signed(-{in[1195-:4],1'b0})+$signed(-{in[1143-:4],1'b0})+$signed(-in[615-:4]);
assign sharing166 = $signed(in[811-:4])+$signed(in[907-:4])+$signed(-{in[1155-:4],1'b0})+$signed(-in[1515-:4])+$signed(-in[471-:4]);
assign sharing167 = $signed(in[1927-:4])+$signed(-{in[1139-:4],1'b0})+$signed(-in[211-:4])+$signed(-in[1231-:4])+$signed(-in[407-:4]);
assign sharing168 = $signed({in[203-:4],1'b0})+$signed(in[111-:4])+$signed(-{in[1539-:4],1'b0})+$signed(-in[1323-:4])+$signed(-in[1683-:4])+$signed(-{in[1591-:4],1'b0})+$signed(-{in[1535-:4],2'b0});
assign sharing169 = $signed(in[1651-:4])+$signed(in[675-:4])+$signed(in[2007-:4])+$signed(-in[1059-:4])+$signed(-in[1619-:4])+$signed(-in[523-:4]);
assign sharing170 = $signed(in[1959-:4])+$signed(in[1135-:4])+$signed({in[415-:4],1'b0})+$signed(in[1055-:4]);
assign sharing171 = $signed(in[1751-:4])+$signed(in[87-:4])+$signed(-in[267-:4]);
assign sharing172 = $signed(in[619-:4])+$signed(in[1699-:4])+$signed({in[815-:4],1'b0})+$signed(in[807-:4])+$signed(-{in[355-:4],1'b0})+$signed(-in[1683-:4])+$signed(-in[327-:4]);
assign sharing173 = $signed(in[1075-:4])+$signed(in[819-:4])+$signed(in[1155-:4])+$signed(in[499-:4])+$signed(-in[471-:4]);
assign sharing174 = $signed({in[1611-:4],1'b0})+$signed(in[1799-:4])+$signed(in[1167-:4]);
assign sharing175 = $signed({in[1675-:4],2'b0})+$signed(in[943-:4])+$signed(-in[387-:4])+$signed(-in[1831-:4]);
assign sharing176 = $signed({in[971-:4],1'b0})+$signed(-{in[91-:4],1'b0})+$signed(-{in[1607-:4],1'b0})+$signed(-in[87-:4]);
assign sharing177 = $signed(in[1547-:4])+$signed(-in[175-:4])+$signed(-in[555-:4])+$signed(-{in[1519-:4],1'b0})+$signed(-in[215-:4]);
assign sharing178 = $signed({in[1827-:4],1'b0})+$signed({in[527-:4],1'b0})+$signed(-in[571-:4]);
assign sharing179 = $signed(in[1967-:4])+$signed(in[603-:4])+$signed(in[655-:4])+$signed(-in[1011-:4]);
assign sharing180 = $signed({in[1483-:4],1'b0})+$signed({in[947-:4],1'b0})+$signed({in[1587-:4],1'b0})+$signed(-in[43-:4])+$signed(-in[911-:4]);
assign sharing181 = $signed(in[1067-:4])+$signed(in[1507-:4])+$signed(in[1031-:4]);
assign sharing182 = $signed({in[1739-:4],1'b0})+$signed(in[119-:4])+$signed({in[1751-:4],1'b0})+$signed(in[407-:4])+$signed(in[1631-:4])+$signed(-{in[2019-:4],1'b0})+$signed(-in[1351-:4]);
assign sharing183 = $signed(in[1539-:4])+$signed(in[1171-:4])+$signed(in[1847-:4])+$signed(-{in[75-:4],2'b0})+$signed(-{in[799-:4],1'b0});
assign sharing184 = $signed({in[1723-:4],1'b0})+$signed(in[995-:4])+$signed(in[319-:4])+$signed(-in[1287-:4]);
assign sharing185 = $signed(in[643-:4])+$signed(in[1383-:4])+$signed(-in[1247-:4]);
assign sharing186 = $signed(in[967-:4])+$signed(in[1903-:4])+$signed(-in[299-:4])+$signed(-{in[1343-:4],1'b0})+$signed(-in[615-:4]);
assign sharing187 = $signed({in[1763-:4],1'b0})+$signed(in[215-:4])+$signed(-in[191-:4]);
assign sharing188 = $signed({in[1875-:4],1'b0})+$signed(in[1331-:4])+$signed({in[1919-:4],1'b0})+$signed(in[2027-:4]);
assign sharing189 = $signed(in[323-:4])+$signed(in[1219-:4])+$signed(-in[115-:4])+$signed(-{in[1735-:4],2'b0});
assign sharing190 = $signed({in[759-:4],1'b0})+$signed(-in[287-:4])+$signed(-in[223-:4]);
assign sharing191 = $signed({in[1419-:4],1'b0})+$signed(in[811-:4])+$signed({in[1431-:4],1'b0})+$signed(in[491-:4])+$signed(-{in[635-:4],1'b0});
assign sharing192 = $signed(in[311-:4])+$signed(-{in[1123-:4],1'b0})+$signed(-in[751-:4])+$signed(-{in[1127-:4],1'b0})+$signed(-in[159-:4]);
assign sharing193 = $signed(in[507-:4])+$signed({in[1503-:4],1'b0})+$signed(-in[291-:4])+$signed(-{in[1671-:4],1'b0})+$signed(-in[423-:4]);
assign sharing194 = $signed(in[391-:4])+$signed(in[915-:4])+$signed(in[863-:4])+$signed(in[1711-:4])+$signed(-in[659-:4])+$signed(-in[271-:4]);
assign sharing195 = $signed(-in[1051-:4])+$signed(-in[907-:4])+$signed(-in[375-:4]);
assign sharing196 = $signed(in[823-:4])+$signed({in[1887-:4],1'b0})+$signed(in[535-:4]);
assign sharing197 = $signed({in[1847-:4],1'b0})+$signed(-in[1747-:4])+$signed(-in[359-:4]);
assign sharing198 = $signed(in[1387-:4])+$signed(in[1347-:4])+$signed(in[259-:4])+$signed(in[1735-:4])+$signed(-in[247-:4]);
assign sharing199 = $signed(in[503-:4])+$signed(-in[851-:4])+$signed(-in[195-:4])+$signed(-in[1503-:4]);
assign sharing200 = $signed(in[951-:4])+$signed(in[1703-:4])+$signed(-in[479-:4]);
assign sharing201 = $signed(in[963-:4])+$signed({in[619-:4],1'b0})+$signed({in[1295-:4],1'b0})+$signed({in[1299-:4],1'b0})+$signed({in[567-:4],1'b0})+$signed(-in[307-:4])+$signed(-in[1455-:4]);
assign sharing202 = $signed({in[1039-:4],1'b0})+$signed({in[1439-:4],1'b0})+$signed(in[103-:4])+$signed(-in[799-:4]);
assign sharing203 = $signed(in[895-:4])+$signed(-in[1159-:4])+$signed(-in[1087-:4])+$signed(-in[463-:4]);
assign sharing204 = $signed(in[315-:4])+$signed(in[311-:4])+$signed({in[1983-:4],1'b0})+$signed(in[255-:4])+$signed(-{in[83-:4],2'b0})+$signed(-in[755-:4]);
assign sharing205 = $signed(in[35-:4])+$signed(-in[443-:4])+$signed(-{in[2015-:4],1'b0});
assign sharing206 = $signed({in[955-:4],1'b0})+$signed(in[243-:4])+$signed(in[775-:4])+$signed(in[1275-:4])+$signed(-{in[259-:4],1'b0})+$signed(-in[1427-:4]);
assign sharing207 = $signed(in[659-:4])+$signed(-in[1783-:4])+$signed(-in[367-:4]);
assign sharing208 = $signed(in[39-:4])+$signed(-{in[459-:4],1'b0})+$signed(-in[1803-:4]);
assign sharing209 = $signed(in[531-:4])+$signed(in[1971-:4])+$signed({in[1559-:4],1'b0})+$signed(-in[1019-:4]);
assign sharing210 = $signed(in[527-:4])+$signed(in[1943-:4])+$signed(-{in[1835-:4],1'b0})+$signed(-in[851-:4])+$signed(-in[1435-:4])+$signed(-in[1491-:4]);
assign sharing211 = $signed(in[1107-:4])+$signed(in[1615-:4])+$signed(-in[1183-:4])+$signed(-in[1143-:4]);
assign sharing212 = $signed({in[1215-:4],1'b0})+$signed({in[639-:4],1'b0})+$signed(-in[1675-:4]);
assign sharing213 = $signed(in[347-:4])+$signed(-in[323-:4])+$signed(-in[1055-:4]);
assign sharing214 = $signed({in[1003-:4],1'b0})+$signed(in[1227-:4])+$signed(in[999-:4])+$signed(-in[1915-:4]);
assign sharing215 = $signed(in[1559-:4])+$signed(-{in[299-:4],1'b0})+$signed(-in[1483-:4])+$signed(-in[1255-:4]);
assign sharing216 = $signed(in[1811-:4])+$signed(-in[1151-:4])+$signed(-in[359-:4]);
assign sharing217 = $signed({in[1347-:4],1'b0})+$signed(in[2011-:4])+$signed({in[1159-:4],1'b0})+$signed({in[255-:4],1'b0})+$signed(-in[851-:4])+$signed(-in[467-:4]);
assign sharing218 = $signed({in[923-:4],1'b0})+$signed({in[1991-:4],1'b0})+$signed(in[591-:4])+$signed(-{in[1819-:4],2'b0})+$signed(-{in[519-:4],2'b0})+$signed(-{in[415-:4],2'b0});
assign sharing219 = $signed({in[1671-:4],1'b0})+$signed(-{in[1955-:4],1'b0})+$signed(-{in[1491-:4],1'b0})+$signed(-{in[1951-:4],1'b0});
assign sharing220 = $signed({in[811-:4],1'b0})+$signed(in[1863-:4])+$signed(in[1279-:4])+$signed(-{in[1883-:4],1'b0});
assign sharing221 = $signed(in[1839-:4])+$signed(in[1567-:4])+$signed(-{in[1567-:4],2'b0});
assign sharing222 = $signed({in[203-:4],2'b0})+$signed(in[1779-:4])+$signed(in[1015-:4]);
assign sharing223 = $signed(in[1819-:4])+$signed(in[151-:4])+$signed(-{in[1819-:4],2'b0})+$signed(-{in[1055-:4],2'b0});
assign sharing224 = $signed({in[459-:4],1'b0})+$signed(-in[75-:4])+$signed(-in[1755-:4]);
assign sharing225 = $signed(in[819-:4])+$signed(in[1135-:4])+$signed(in[327-:4])+$signed(-in[655-:4]);
assign sharing226 = $signed({in[475-:4],1'b0})+$signed(in[1311-:4])+$signed(-{in[259-:4],2'b0});
assign sharing227 = $signed(in[131-:4])+$signed(in[2019-:4])+$signed(-in[903-:4]);
assign sharing228 = $signed(in[1091-:4])+$signed(in[1331-:4])+$signed(in[1007-:4])+$signed(-in[531-:4])+$signed(-in[295-:4]);
assign sharing229 = $signed(in[1879-:4])+$signed({in[1975-:4],1'b0})+$signed(in[239-:4])+$signed(-{in[1463-:4],1'b0});
assign sharing230 = $signed(in[147-:4])+$signed(-in[1227-:4])+$signed(-in[1655-:4]);
assign sharing231 = $signed(in[1179-:4])+$signed(in[1715-:4])+$signed(in[1235-:4])+$signed(-in[103-:4]);
assign sharing232 = $signed({in[267-:4],1'b0})+$signed({in[999-:4],1'b0})+$signed(-in[1975-:4]);
assign sharing233 = $signed(-{in[1059-:4],1'b0})+$signed(-{in[1091-:4],1'b0})+$signed(-{in[1863-:4],1'b0})+$signed(-{in[1615-:4],2'b0})+$signed(-{in[1107-:4],2'b0});
assign sharing234 = $signed({in[867-:4],1'b0})+$signed(in[947-:4])+$signed(in[79-:4])+$signed(-{in[1595-:4],1'b0})+$signed(-{in[1599-:4],1'b0});
assign sharing235 = $signed(in[411-:4])+$signed(in[767-:4])+$signed(-{in[1819-:4],1'b0})+$signed(-in[1495-:4]);
assign sharing236 = $signed({in[1643-:4],1'b0})+$signed({in[1775-:4],1'b0})+$signed(in[1951-:4]);
assign sharing237 = $signed(in[1867-:4])+$signed({in[1487-:4],1'b0})+$signed(in[1439-:4]);
assign sharing238 = $signed(in[1687-:4])+$signed(in[1283-:4])+$signed(in[383-:4])+$signed(-{in[947-:4],1'b0});
assign sharing239 = $signed(in[859-:4])+$signed(-in[1335-:4])+$signed(-in[247-:4]);
assign sharing240 = $signed(in[1607-:4])+$signed(in[1191-:4])+$signed(-in[371-:4]);
assign sharing241 = $signed({in[1595-:4],2'b0})+$signed(-{in[803-:4],1'b0})+$signed(-in[843-:4]);
assign sharing242 = $signed(in[1943-:4])+$signed(in[1643-:4])+$signed(in[883-:4])+$signed(in[223-:4]);
assign sharing243 = $signed(-{in[123-:4],2'b0})+$signed(-in[1931-:4])+$signed(-{in[811-:4],2'b0});
assign sharing244 = $signed(in[1543-:4])+$signed({in[1711-:4],1'b0})+$signed(in[935-:4]);
assign sharing245 = $signed(in[1527-:4])+$signed({in[1207-:4],1'b0})+$signed(in[447-:4]);
assign sharing246 = $signed({in[1291-:4],1'b0})+$signed(in[555-:4])+$signed({in[615-:4],1'b0})+$signed(-in[1519-:4]);
assign sharing247 = $signed({in[443-:4],2'b0})+$signed({in[1843-:4],1'b0})+$signed(in[1871-:4])+$signed(-{in[1515-:4],1'b0});
assign sharing248 = $signed(in[803-:4])+$signed(in[203-:4])+$signed(-in[1815-:4]);
assign sharing249 = $signed({in[1795-:4],1'b0})+$signed(-in[307-:4])+$signed(-in[263-:4]);
assign sharing250 = $signed({in[335-:4],1'b0})+$signed(-in[1239-:4])+$signed(-in[319-:4]);
assign sharing251 = $signed({in[763-:4],1'b0})+$signed({in[771-:4],1'b0})+$signed(in[15-:4])+$signed(-in[1723-:4]);
assign sharing252 = $signed({in[559-:4],1'b0})+$signed({in[1167-:4],1'b0})+$signed({in[135-:4],1'b0})+$signed(in[511-:4]);
assign sharing253 = $signed(in[1647-:4])+$signed(in[751-:4])+$signed(-in[219-:4])+$signed(-in[1267-:4]);
assign sharing254 = $signed({in[483-:4],1'b0})+$signed({in[491-:4],1'b0})+$signed(in[647-:4]);
assign sharing255 = $signed(in[1451-:4])+$signed(-in[283-:4])+$signed(-in[115-:4]);
assign weighted_sum[0] = $signed(-{in[771-:4],2'b0})+$signed(-{in[775-:4],1'b0})+$signed(-in[391-:4])+$signed({in[1803-:4],1'b0})+$signed(in[139-:4])+$signed({in[275-:4],1'b0})+$signed({in[1683-:4],1'b0})+$signed({in[279-:4],1'b0})+$signed(in[151-:4])+$signed({in[1687-:4],1'b0})+$signed(in[1439-:4])+$signed({in[931-:4],1'b0})+$signed(-{in[1443-:4],1'b0})+$signed(-in[1699-:4])+$signed(-{in[1447-:4],1'b0})+$signed(-{in[1451-:4],1'b0})+$signed(-in[1707-:4])+$signed({in[1967-:4],1'b0})+$signed(in[567-:4])+$signed(in[571-:4])+$signed(-{in[1471-:4],2'b0})+$signed({in[1727-:4],1'b0})+$signed(in[1215-:4])+$signed({in[1731-:4],1'b0})+$signed({in[203-:4],1'b0})+$signed(-{in[83-:4],1'b0})+$signed(-in[211-:4])+$signed(-{in[87-:4],1'b0})+$signed({in[1495-:4],1'b0})+$signed({in[1623-:4],1'b0})+$signed({in[1499-:4],1'b0})+$signed(in[859-:4])+$signed({in[1631-:4],1'b0})+$signed(in[607-:4])+$signed(in[1503-:4])+$signed(-{in[99-:4],1'b0})+$signed(-in[1379-:4])+$signed({in[1639-:4],1'b0})+$signed(-in[359-:4])+$signed({in[623-:4],1'b0})+$signed({in[879-:4],1'b0})+$signed(-{in[115-:4],2'b0})+$signed({in[371-:4],1'b0})+$signed(-{in[1523-:4],1'b0})+$signed(-{in[119-:4],1'b0})+$signed(-{in[123-:4],1'b0})+$signed(-{in[895-:4],1'b0})+$signed(sharing0)+$signed(sharing1)+$signed(sharing32)+$signed(sharing33)+$signed(sharing64)+$signed(sharing65)+$signed(sharing96)+$signed(sharing97)+$signed(sharing127)+$signed(sharing128)+$signed(sharing155)+$signed(sharing177)+$signed(sharing201)+$signed(sharing217)+$signed(sharing230)+$signed(sharing236)+$signed(sharing241)+$signed(1);
assign weighted_sum[1] = $signed(in[1923-:4])+$signed(-{in[263-:4],2'b0})+$signed({in[519-:4],1'b0})+$signed(in[1675-:4])+$signed({in[1423-:4],1'b0})+$signed(-{in[403-:4],1'b0})+$signed(-in[1811-:4])+$signed(in[1939-:4])+$signed(in[1947-:4])+$signed(in[27-:4])+$signed(in[155-:4])+$signed(-{in[1695-:4],1'b0})+$signed(in[547-:4])+$signed(-in[1315-:4])+$signed(-{in[1063-:4],1'b0})+$signed({in[555-:4],1'b0})+$signed(in[1583-:4])+$signed(-in[1075-:4])+$signed(in[183-:4])+$signed(-{in[1723-:4],2'b0})+$signed(in[187-:4])+$signed({in[579-:4],1'b0})+$signed({in[1235-:4],1'b0})+$signed(in[595-:4])+$signed(-in[215-:4])+$signed(in[1239-:4])+$signed(-in[1119-:4])+$signed(-in[223-:4])+$signed(in[1503-:4])+$signed(-{in[1507-:4],1'b0})+$signed(in[1635-:4])+$signed({in[359-:4],1'b0})+$signed(-in[1015-:4])+$signed(in[507-:4])+$signed(sharing2)+$signed(sharing3)+$signed(sharing34)+$signed(sharing35)+$signed(sharing66)+$signed(sharing67)+$signed(sharing104)+$signed(-sharing105)+$signed(sharing129)+$signed(sharing130)+$signed(-sharing165)+$signed(sharing178)+$signed(sharing179)+$signed(sharing202)+$signed(-2);
assign weighted_sum[2] = $signed(in[515-:4])+$signed(in[1923-:4])+$signed(-{in[1675-:4],3'b0})+$signed({in[1675-:4],1'b0})+$signed(in[651-:4])+$signed(-{in[271-:4],2'b0})+$signed(-{in[1551-:4],1'b0})+$signed(-{in[275-:4],3'b0})+$signed(-{in[1555-:4],3'b0})+$signed(-{in[279-:4],3'b0})+$signed(-{in[151-:4],1'b0})+$signed(in[1431-:4])+$signed({in[279-:4],1'b0})+$signed(-in[667-:4])+$signed(in[1823-:4])+$signed(in[927-:4])+$signed({in[163-:4],1'b0})+$signed(in[419-:4])+$signed({in[167-:4],1'b0})+$signed(-in[1447-:4])+$signed({in[1579-:4],1'b0})+$signed(in[171-:4])+$signed(-{in[955-:4],2'b0})+$signed(in[187-:4])+$signed(-{in[959-:4],3'b0})+$signed(-{in[319-:4],1'b0})+$signed(-in[703-:4])+$signed({in[1471-:4],1'b0})+$signed(-{in[323-:4],2'b0})+$signed(-in[1727-:4])+$signed(in[1871-:4])+$signed({in[467-:4],1'b0})+$signed(-in[1623-:4])+$signed(-{in[1627-:4],2'b0})+$signed(-{in[987-:4],1'b0})+$signed(-in[1115-:4])+$signed(-{in[1631-:4],3'b0})+$signed(-{in[1503-:4],2'b0})+$signed(-{in[1635-:4],3'b0})+$signed(-{in[227-:4],1'b0})+$signed({in[1635-:4],1'b0})+$signed(-{in[231-:4],1'b0})+$signed(-{in[359-:4],1'b0})+$signed({in[1771-:4],1'b0})+$signed(-in[747-:4])+$signed(-{in[751-:4],1'b0})+$signed(in[247-:4])+$signed({in[635-:4],1'b0})+$signed(in[379-:4])+$signed(in[511-:4])+$signed(sharing24)+$signed(-sharing25)+$signed(sharing36)+$signed(sharing37)+$signed(sharing68)+$signed(sharing69)+$signed(sharing98)+$signed(sharing99)+$signed(-sharing155)+$signed(sharing180)+$signed(sharing226)+$signed(-sharing235)+$signed(sharing237)+$signed(0);
assign weighted_sum[3] = $signed(-in[1923-:4])+$signed({in[1543-:4],1'b0})+$signed(in[519-:4])+$signed(-in[7-:4])+$signed({in[907-:4],1'b0})+$signed(-in[779-:4])+$signed({in[911-:4],1'b0})+$signed(in[271-:4])+$signed({in[403-:4],1'b0})+$signed(-in[19-:4])+$signed({in[531-:4],1'b0})+$signed({in[1555-:4],1'b0})+$signed(in[1683-:4])+$signed(-in[1435-:4])+$signed({in[1699-:4],1'b0})+$signed(-in[675-:4])+$signed(in[1831-:4])+$signed(-in[1959-:4])+$signed({in[299-:4],1'b0})+$signed(in[939-:4])+$signed(-{in[1195-:4],1'b0})+$signed(in[1711-:4])+$signed({in[1595-:4],1'b0})+$signed(-in[443-:4])+$signed({in[831-:4],1'b0})+$signed(in[1727-:4])+$signed({in[323-:4],1'b0})+$signed({in[1603-:4],1'b0})+$signed({in[1735-:4],1'b0})+$signed(in[583-:4])+$signed({in[587-:4],1'b0})+$signed({in[1611-:4],1'b0})+$signed(-{in[1867-:4],1'b0})+$signed(-{in[1871-:4],2'b0})+$signed(-{in[79-:4],1'b0})+$signed({in[975-:4],1'b0})+$signed(-{in[467-:4],2'b0})+$signed(-in[1107-:4])+$signed({in[987-:4],1'b0})+$signed(in[759-:4])+$signed(-in[627-:4])+$signed(-{in[759-:4],2'b0})+$signed(-{in[1143-:4],1'b0})+$signed(in[247-:4])+$signed(-in[1023-:4])+$signed(sharing4)+$signed(sharing5)+$signed(sharing32)+$signed(-sharing33)+$signed(sharing72)+$signed(-sharing73)+$signed(sharing100)+$signed(sharing101)+$signed(sharing131)+$signed(sharing164)+$signed(sharing181)+$signed(sharing182)+$signed(sharing203)+$signed(sharing218)+$signed(sharing231)+$signed(sharing242)+$signed(sharing248)+$signed(1);
assign weighted_sum[4] = $signed(-{in[515-:4],2'b0})+$signed(in[1543-:4])+$signed({in[639-:4],1'b0})+$signed(-{in[1423-:4],1'b0})+$signed({in[659-:4],2'b0})+$signed(in[1947-:4])+$signed(-in[539-:4])+$signed(in[1567-:4])+$signed(in[931-:4])+$signed(in[1955-:4])+$signed(-in[1447-:4])+$signed(in[1575-:4])+$signed({in[1323-:4],1'b0})+$signed(-in[1451-:4])+$signed({in[1327-:4],1'b0})+$signed({in[1331-:4],2'b0})+$signed(-{in[1207-:4],1'b0})+$signed(in[183-:4])+$signed(-{in[571-:4],1'b0})+$signed(-in[1467-:4])+$signed(-{in[67-:4],2'b0})+$signed(in[579-:4])+$signed({in[1995-:4],1'b0})+$signed({in[1999-:4],1'b0})+$signed(-{in[467-:4],1'b0})+$signed(in[1491-:4])+$signed({in[2003-:4],1'b0})+$signed(-{in[87-:4],2'b0})+$signed(-{in[91-:4],2'b0})+$signed({in[603-:4],1'b0})+$signed(in[1115-:4])+$signed({in[2011-:4],2'b0})+$signed(-{in[479-:4],1'b0})+$signed(in[871-:4])+$signed(in[235-:4])+$signed(-in[1515-:4])+$signed(in[1519-:4])+$signed(-in[1775-:4])+$signed(-{in[1911-:4],1'b0})+$signed({in[1531-:4],1'b0})+$signed(in[1787-:4])+$signed(-{in[1919-:4],1'b0})+$signed(sharing0)+$signed(-sharing1)+$signed(sharing38)+$signed(sharing39)+$signed(sharing92)+$signed(-sharing93)+$signed(sharing102)+$signed(sharing103)+$signed(sharing132)+$signed(sharing133)+$signed(sharing161)+$signed(-sharing191)+$signed(sharing204)+$signed(sharing218)+$signed(sharing238)+$signed(1);
assign weighted_sum[5] = $signed({in[771-:4],1'b0})+$signed(-in[1927-:4])+$signed(-in[135-:4])+$signed(in[395-:4])+$signed(-{in[1935-:4],2'b0})+$signed(-{in[1939-:4],1'b0})+$signed(-in[531-:4])+$signed(in[1171-:4])+$signed(in[1299-:4])+$signed(in[1559-:4])+$signed(-in[1687-:4])+$signed(in[151-:4])+$signed(-in[291-:4])+$signed(in[1315-:4])+$signed(-in[1827-:4])+$signed(-{in[1575-:4],1'b0})+$signed(-in[1955-:4])+$signed(-{in[1579-:4],2'b0})+$signed(in[1835-:4])+$signed(-in[1071-:4])+$signed(-{in[311-:4],2'b0})+$signed({in[959-:4],1'b0})+$signed(-in[1475-:4])+$signed(in[331-:4])+$signed(-in[975-:4])+$signed(in[1743-:4])+$signed(-{in[599-:4],1'b0})+$signed(-{in[987-:4],2'b0})+$signed(in[347-:4])+$signed(-in[1499-:4])+$signed(-{in[223-:4],1'b0})+$signed({in[2023-:4],1'b0})+$signed(in[1127-:4])+$signed(-in[1003-:4])+$signed(-{in[1647-:4],2'b0})+$signed(-{in[1651-:4],2'b0})+$signed(-{in[1527-:4],1'b0})+$signed(in[631-:4])+$signed({in[1783-:4],1'b0})+$signed(-{in[1531-:4],1'b0})+$signed(-in[1019-:4])+$signed(-{in[1663-:4],2'b0})+$signed(-{in[895-:4],1'b0})+$signed(sharing4)+$signed(-sharing5)+$signed(sharing54)+$signed(-sharing55)+$signed(sharing70)+$signed(sharing71)+$signed(sharing106)+$signed(-sharing107)+$signed(sharing145)+$signed(-sharing146)+$signed(sharing156)+$signed(sharing157)+$signed(-sharing180)+$signed(-sharing232)+$signed(-sharing236)+$signed(-sharing255)+$signed(2);
assign weighted_sum[6] = $signed(-{in[387-:4],2'b0})+$signed({in[1667-:4],1'b0})+$signed(-in[1795-:4])+$signed(-{in[383-:4],1'b0})+$signed(-in[1543-:4])+$signed(in[1287-:4])+$signed(-in[395-:4])+$signed(-in[143-:4])+$signed(-in[1039-:4])+$signed(in[1679-:4])+$signed(-{in[1427-:4],1'b0})+$signed(in[275-:4])+$signed(-in[403-:4])+$signed({in[1811-:4],1'b0})+$signed(in[1563-:4])+$signed(-in[1691-:4])+$signed({in[287-:4],1'b0})+$signed(-{in[1831-:4],1'b0})+$signed(in[167-:4])+$signed(-{in[1067-:4],3'b0})+$signed(-{in[427-:4],2'b0})+$signed({in[1067-:4],1'b0})+$signed(-{in[431-:4],2'b0})+$signed(-{in[1839-:4],1'b0})+$signed(-{in[435-:4],1'b0})+$signed(-in[1847-:4])+$signed(-in[1851-:4])+$signed(in[959-:4])+$signed(-{in[1743-:4],3'b0})+$signed(-{in[79-:4],1'b0})+$signed(in[1103-:4])+$signed(-{in[339-:4],2'b0})+$signed(-in[1879-:4])+$signed({in[219-:4],1'b0})+$signed(-{in[1115-:4],1'b0})+$signed(-in[1243-:4])+$signed(-{in[1119-:4],2'b0})+$signed({in[223-:4],1'b0})+$signed(-in[863-:4])+$signed(-in[483-:4])+$signed(in[1259-:4])+$signed(-{in[1779-:4],1'b0})+$signed(-in[1019-:4])+$signed(-{in[1791-:4],2'b0})+$signed(-{in[895-:4],1'b0})+$signed(sharing12)+$signed(-sharing13)+$signed(sharing60)+$signed(-sharing61)+$signed(sharing78)+$signed(-sharing79)+$signed(sharing98)+$signed(-sharing99)+$signed(sharing153)+$signed(-sharing154)+$signed(sharing170)+$signed(-sharing171)+$signed(-sharing177)+$signed(sharing210)+$signed(sharing220)+$signed(-sharing248)+$signed(2);
assign weighted_sum[7] = $signed(in[387-:4])+$signed(-{in[1163-:4],2'b0})+$signed(-{in[1035-:4],1'b0})+$signed(in[267-:4])+$signed(-{in[1167-:4],2'b0})+$signed(in[1043-:4])+$signed(in[1171-:4])+$signed(-{in[1175-:4],2'b0})+$signed(in[1307-:4])+$signed(in[1823-:4])+$signed(-{in[1831-:4],2'b0})+$signed(-in[423-:4])+$signed(-{in[1835-:4],2'b0})+$signed(in[1323-:4])+$signed(in[1707-:4])+$signed(-{in[1839-:4],1'b0})+$signed(-{in[307-:4],1'b0})+$signed(-in[435-:4])+$signed(in[1331-:4])+$signed(in[567-:4])+$signed(-in[1079-:4])+$signed(in[1595-:4])+$signed(-{in[1215-:4],3'b0})+$signed({in[1727-:4],1'b0})+$signed(-{in[1219-:4],3'b0})+$signed({in[1219-:4],1'b0})+$signed(in[1731-:4])+$signed(-{in[1223-:4],2'b0})+$signed(in[1231-:4])+$signed(in[2003-:4])+$signed(in[599-:4])+$signed(-in[983-:4])+$signed(-in[987-:4])+$signed(in[1499-:4])+$signed(-{in[479-:4],2'b0})+$signed(-{in[483-:4],3'b0})+$signed(-{in[487-:4],3'b0})+$signed(-{in[1895-:4],2'b0})+$signed(in[999-:4])+$signed(-{in[491-:4],3'b0})+$signed(-{in[1899-:4],2'b0})+$signed(in[1899-:4])+$signed(-{in[495-:4],2'b0})+$signed({in[1263-:4],1'b0})+$signed(in[623-:4])+$signed(in[379-:4])+$signed({in[1791-:4],1'b0})+$signed(sharing18)+$signed(-sharing19)+$signed(sharing48)+$signed(-sharing49)+$signed(sharing82)+$signed(-sharing83)+$signed(sharing100)+$signed(-sharing101)+$signed(sharing134)+$signed(-sharing135)+$signed(-sharing173)+$signed(sharing192)+$signed(sharing212)+$signed(-sharing213)+$signed(sharing254)+$signed(2);
assign weighted_sum[8] = $signed(-{in[131-:4],3'b0})+$signed(in[131-:4])+$signed(-{in[135-:4],3'b0})+$signed(in[1527-:4])+$signed(-{in[139-:4],2'b0})+$signed({in[651-:4],1'b0})+$signed(-in[1291-:4])+$signed(-{in[143-:4],2'b0})+$signed(-{in[1935-:4],2'b0})+$signed(-{in[1939-:4],2'b0})+$signed(-{in[535-:4],2'b0})+$signed(-{in[1943-:4],2'b0})+$signed(-{in[539-:4],1'b0})+$signed(-{in[1947-:4],1'b0})+$signed(in[671-:4])+$signed(-{in[803-:4],2'b0})+$signed(in[1059-:4])+$signed(-{in[807-:4],2'b0})+$signed(-{in[815-:4],2'b0})+$signed(-in[559-:4])+$signed(-{in[819-:4],2'b0})+$signed(in[179-:4])+$signed(-{in[823-:4],1'b0})+$signed(in[1719-:4])+$signed(-{in[1467-:4],1'b0})+$signed(-{in[1471-:4],2'b0})+$signed({in[319-:4],1'b0})+$signed(-{in[1475-:4],2'b0})+$signed(-{in[71-:4],2'b0})+$signed(-{in[1479-:4],2'b0})+$signed(in[1991-:4])+$signed(-{in[1483-:4],2'b0})+$signed(-{in[79-:4],2'b0})+$signed(-{in[1487-:4],2'b0})+$signed(in[79-:4])+$signed(in[1747-:4])+$signed(-{in[855-:4],2'b0})+$signed(-{in[91-:4],1'b0})+$signed(-in[1499-:4])+$signed(-in[2015-:4])+$signed(-{in[1907-:4],1'b0})+$signed(-{in[119-:4],1'b0})+$signed(in[1783-:4])+$signed(in[1531-:4])+$signed(-{in[127-:4],3'b0})+$signed({in[1535-:4],1'b0})+$signed(in[127-:4])+$signed(sharing6)+$signed(sharing7)+$signed(sharing40)+$signed(sharing41)+$signed(sharing72)+$signed(sharing73)+$signed(sharing104)+$signed(sharing105)+$signed(sharing139)+$signed(-sharing140)+$signed(sharing158)+$signed(sharing183)+$signed(sharing184)+$signed(sharing204)+$signed(sharing219)+$signed(sharing232)+$signed(sharing243)+$signed(2);
assign weighted_sum[9] = $signed(-in[1671-:4])+$signed(in[779-:4])+$signed({in[1423-:4],1'b0})+$signed(-in[1167-:4])+$signed(in[527-:4])+$signed({in[1427-:4],1'b0})+$signed(-in[1811-:4])+$signed({in[1431-:4],1'b0})+$signed(in[1943-:4])+$signed(in[407-:4])+$signed({in[1435-:4],1'b0})+$signed({in[539-:4],1'b0})+$signed(-in[419-:4])+$signed(in[1703-:4])+$signed({in[1579-:4],1'b0})+$signed(in[171-:4])+$signed(-in[427-:4])+$signed(-in[431-:4])+$signed(in[951-:4])+$signed(in[1591-:4])+$signed(-in[1847-:4])+$signed(in[703-:4])+$signed({in[67-:4],1'b0})+$signed({in[71-:4],1'b0})+$signed(-{in[327-:4],1'b0})+$signed(in[75-:4])+$signed(in[459-:4])+$signed({in[1871-:4],1'b0})+$signed(-in[1103-:4])+$signed({in[1887-:4],1'b0})+$signed(-in[1119-:4])+$signed({in[1895-:4],1'b0})+$signed(in[103-:4])+$signed(-in[871-:4])+$signed({in[363-:4],1'b0})+$signed(in[1131-:4])+$signed({in[1899-:4],1'b0})+$signed(-in[879-:4])+$signed({in[1143-:4],1'b0})+$signed(sharing8)+$signed(sharing9)+$signed(sharing42)+$signed(sharing43)+$signed(sharing74)+$signed(sharing75)+$signed(sharing106)+$signed(sharing107)+$signed(sharing134)+$signed(sharing135)+$signed(sharing159)+$signed(sharing160)+$signed(sharing185)+$signed(sharing186)+$signed(sharing205)+$signed(-sharing217)+$signed(1);
assign weighted_sum[10] = $signed({in[515-:4],1'b0})+$signed(in[1923-:4])+$signed({in[519-:4],1'b0})+$signed(in[907-:4])+$signed(in[403-:4])+$signed(-in[531-:4])+$signed(-in[1939-:4])+$signed({in[1819-:4],1'b0})+$signed(in[1951-:4])+$signed(-in[31-:4])+$signed(in[799-:4])+$signed(in[1955-:4])+$signed({in[807-:4],1'b0})+$signed(-in[935-:4])+$signed({in[171-:4],1'b0})+$signed({in[815-:4],1'b0})+$signed({in[439-:4],1'b0})+$signed(in[439-:4])+$signed(in[823-:4])+$signed({in[1479-:4],1'b0})+$signed(in[459-:4])+$signed({in[1871-:4],1'b0})+$signed(in[2003-:4])+$signed({in[855-:4],1'b0})+$signed(in[599-:4])+$signed({in[2007-:4],1'b0})+$signed({in[95-:4],1'b0})+$signed({in[1119-:4],1'b0})+$signed(in[1247-:4])+$signed(in[99-:4])+$signed(-in[235-:4])+$signed(in[875-:4])+$signed(in[883-:4])+$signed(in[1523-:4])+$signed(in[759-:4])+$signed(in[1531-:4])+$signed(sharing10)+$signed(sharing11)+$signed(sharing44)+$signed(sharing45)+$signed(sharing76)+$signed(sharing77)+$signed(sharing108)+$signed(sharing109)+$signed(sharing136)+$signed(sharing137)+$signed(-sharing158)+$signed(sharing187)+$signed(sharing188)+$signed(-sharing205)+$signed(sharing220)+$signed(sharing234)+$signed(sharing252)+$signed(0);
assign weighted_sum[11] = $signed({in[1923-:4],1'b0})+$signed(in[1667-:4])+$signed({in[267-:4],1'b0})+$signed({in[1039-:4],1'b0})+$signed({in[1295-:4],1'b0})+$signed(-{in[1679-:4],1'b0})+$signed(in[1935-:4])+$signed(-{in[1683-:4],1'b0})+$signed(in[19-:4])+$signed(-{in[1687-:4],2'b0})+$signed(-in[663-:4])+$signed(in[1175-:4])+$signed(-in[1307-:4])+$signed(in[539-:4])+$signed({in[1055-:4],1'b0})+$signed(-in[675-:4])+$signed(in[1319-:4])+$signed(-in[1831-:4])+$signed(in[1839-:4])+$signed(-{in[1715-:4],1'b0})+$signed(in[435-:4])+$signed(-in[1587-:4])+$signed({in[1971-:4],1'b0})+$signed(-in[311-:4])+$signed(in[827-:4])+$signed(-in[1607-:4])+$signed(-{in[1611-:4],2'b0})+$signed(-{in[1743-:4],2'b0})+$signed(-in[207-:4])+$signed({in[211-:4],1'b0})+$signed(in[979-:4])+$signed(-{in[1751-:4],1'b0})+$signed(-{in[475-:4],1'b0})+$signed(-in[219-:4])+$signed(in[1115-:4])+$signed({in[763-:4],1'b0})+$signed(-{in[1639-:4],1'b0})+$signed(in[619-:4])+$signed({in[375-:4],1'b0})+$signed({in[379-:4],1'b0})+$signed(-{in[1663-:4],2'b0})+$signed(sharing12)+$signed(sharing13)+$signed(sharing46)+$signed(sharing47)+$signed(sharing76)+$signed(-sharing77)+$signed(sharing124)+$signed(-sharing125)+$signed(sharing143)+$signed(-sharing144)+$signed(sharing159)+$signed(-sharing160)+$signed(sharing189)+$signed(sharing190)+$signed(sharing206)+$signed(-sharing249)+$signed(2);
assign weighted_sum[12] = $signed(-in[255-:4])+$signed(-in[1927-:4])+$signed(in[903-:4])+$signed(-{in[1555-:4],2'b0})+$signed({in[1815-:4],1'b0})+$signed(in[535-:4])+$signed(in[919-:4])+$signed(-{in[1691-:4],3'b0})+$signed({in[1563-:4],1'b0})+$signed(-{in[1823-:4],2'b0})+$signed(-{in[1055-:4],2'b0})+$signed(-{in[1059-:4],2'b0})+$signed(in[163-:4])+$signed(in[547-:4])+$signed(-in[423-:4])+$signed(-{in[1707-:4],1'b0})+$signed(in[1071-:4])+$signed(in[51-:4])+$signed(-in[823-:4])+$signed(-{in[1723-:4],2'b0})+$signed(in[1723-:4])+$signed(-{in[1727-:4],3'b0})+$signed(in[1215-:4])+$signed(-{in[1731-:4],3'b0})+$signed(in[1983-:4])+$signed({in[1475-:4],1'b0})+$signed(-{in[327-:4],3'b0})+$signed({in[327-:4],1'b0})+$signed(in[1479-:4])+$signed(-{in[331-:4],3'b0})+$signed(-{in[1607-:4],1'b0})+$signed(in[1483-:4])+$signed(-{in[335-:4],3'b0})+$signed(-{in[1103-:4],1'b0})+$signed(in[1615-:4])+$signed(in[467-:4])+$signed(in[1111-:4])+$signed(-in[2015-:4])+$signed(-in[355-:4])+$signed(in[1643-:4])+$signed(-{in[371-:4],2'b0})+$signed(-{in[375-:4],3'b0})+$signed(-{in[1015-:4],2'b0})+$signed(-in[1143-:4])+$signed(-{in[379-:4],2'b0})+$signed(in[1915-:4])+$signed(-in[763-:4])+$signed(in[1535-:4])+$signed(sharing14)+$signed(sharing15)+$signed(sharing36)+$signed(-sharing37)+$signed(sharing78)+$signed(sharing79)+$signed(sharing110)+$signed(sharing111)+$signed(sharing138)+$signed(sharing161)+$signed(sharing189)+$signed(-sharing190)+$signed(sharing216)+$signed(-sharing231)+$signed(sharing245)+$signed(sharing250)+$signed(1);
assign weighted_sum[13] = $signed(-{in[263-:4],1'b0})+$signed(-{in[519-:4],1'b0})+$signed(-{in[1807-:4],2'b0})+$signed({in[911-:4],1'b0})+$signed(-in[143-:4])+$signed(-in[271-:4])+$signed(-{in[147-:4],2'b0})+$signed(-{in[1551-:4],1'b0})+$signed(-in[1427-:4])+$signed(-{in[1555-:4],2'b0})+$signed(-{in[151-:4],2'b0})+$signed(-{in[1811-:4],2'b0})+$signed(-{in[1051-:4],1'b0})+$signed(-in[411-:4])+$signed(-in[155-:4])+$signed(in[1023-:4])+$signed(-{in[1571-:4],2'b0})+$signed(-{in[163-:4],1'b0})+$signed(-{in[167-:4],2'b0})+$signed(-{in[935-:4],2'b0})+$signed(-{in[1575-:4],2'b0})+$signed(-{in[171-:4],2'b0})+$signed({in[1067-:4],1'b0})+$signed(-{in[1711-:4],2'b0})+$signed(-in[943-:4])+$signed(in[187-:4])+$signed(-in[1467-:4])+$signed({in[1599-:4],1'b0})+$signed(-in[831-:4])+$signed(-{in[1859-:4],2'b0})+$signed(-{in[1607-:4],2'b0})+$signed(-{in[1867-:4],2'b0})+$signed(-{in[847-:4],2'b0})+$signed(-in[463-:4])+$signed(-{in[215-:4],2'b0})+$signed(in[343-:4])+$signed({in[859-:4],1'b0})+$signed(in[2015-:4])+$signed(-{in[1763-:4],2'b0})+$signed(-in[611-:4])+$signed(in[2023-:4])+$signed(-{in[875-:4],1'b0})+$signed(-in[107-:4])+$signed(in[491-:4])+$signed(-in[1259-:4])+$signed(-{in[1519-:4],2'b0})+$signed({in[2027-:4],1'b0})+$signed(-{in[1523-:4],3'b0})+$signed(in[1523-:4])+$signed(-{in[1527-:4],3'b0})+$signed({in[1527-:4],1'b0})+$signed(-{in[1659-:4],1'b0})+$signed(in[123-:4])+$signed(-{in[255-:4],2'b0})+$signed(in[1279-:4])+$signed(sharing16)+$signed(sharing17)+$signed(sharing48)+$signed(sharing49)+$signed(sharing86)+$signed(-sharing87)+$signed(sharing126)+$signed(sharing127)+$signed(-sharing128)+$signed(sharing162)+$signed(sharing163)+$signed(sharing185)+$signed(-sharing186)+$signed(sharing207)+$signed(sharing208)+$signed(sharing221)+$signed(-sharing222)+$signed(sharing233)+$signed(-sharing238)+$signed(sharing240)+$signed(sharing243)+$signed(-1);
assign weighted_sum[14] = $signed(-{in[387-:4],1'b0})+$signed(in[259-:4])+$signed(-in[1031-:4])+$signed(in[139-:4])+$signed(-{in[1039-:4],2'b0})+$signed(-in[19-:4])+$signed(in[403-:4])+$signed(-in[23-:4])+$signed(in[1947-:4])+$signed(-in[1563-:4])+$signed(in[671-:4])+$signed(in[163-:4])+$signed(in[931-:4])+$signed(in[1315-:4])+$signed(-{in[307-:4],2'b0})+$signed(-{in[435-:4],2'b0})+$signed(-{in[439-:4],3'b0})+$signed({in[439-:4],1'b0})+$signed(-in[1719-:4])+$signed(in[1475-:4])+$signed(in[1987-:4])+$signed({in[1735-:4],1'b0})+$signed({in[75-:4],1'b0})+$signed(in[1611-:4])+$signed(-{in[1111-:4],3'b0})+$signed(-{in[983-:4],1'b0})+$signed({in[1111-:4],1'b0})+$signed(-{in[1115-:4],3'b0})+$signed(in[119-:4])+$signed(in[91-:4])+$signed(-{in[1119-:4],2'b0})+$signed(-in[1375-:4])+$signed(-{in[1123-:4],2'b0})+$signed(-in[355-:4])+$signed(-{in[359-:4],3'b0})+$signed(in[1507-:4])+$signed({in[359-:4],1'b0})+$signed(in[487-:4])+$signed(-{in[363-:4],1'b0})+$signed(-{in[1783-:4],2'b0})+$signed(-in[1655-:4])+$signed(-{in[1787-:4],2'b0})+$signed(-{in[383-:4],2'b0})+$signed(in[895-:4])+$signed(sharing18)+$signed(sharing19)+$signed(sharing50)+$signed(-sharing51)+$signed(sharing94)+$signed(-sharing95)+$signed(sharing116)+$signed(-sharing117)+$signed(sharing147)+$signed(-sharing148)+$signed(sharing162)+$signed(-sharing163)+$signed(sharing196)+$signed(-sharing197)+$signed(sharing209)+$signed(-sharing247)+$signed(1);
assign weighted_sum[15] = $signed(in[1795-:4])+$signed(-{in[1671-:4],2'b0})+$signed(in[139-:4])+$signed(-{in[659-:4],1'b0})+$signed(-in[915-:4])+$signed(-in[1555-:4])+$signed({in[1687-:4],1'b0})+$signed(-in[919-:4])+$signed(-in[923-:4])+$signed(-in[671-:4])+$signed(-{in[1315-:4],2'b0})+$signed(-{in[1571-:4],1'b0})+$signed(-{in[1955-:4],1'b0})+$signed({in[423-:4],1'b0})+$signed(-{in[1319-:4],1'b0})+$signed(-{in[1323-:4],2'b0})+$signed(-{in[1327-:4],2'b0})+$signed(-in[175-:4])+$signed(in[47-:4])+$signed(-{in[1331-:4],1'b0})+$signed(in[1851-:4])+$signed(-{in[319-:4],2'b0})+$signed(-{in[323-:4],2'b0})+$signed(-{in[1991-:4],2'b0})+$signed(-{in[583-:4],1'b0})+$signed(-in[199-:4])+$signed(in[71-:4])+$signed(-{in[1995-:4],2'b0})+$signed(-{in[1999-:4],2'b0})+$signed(-in[1231-:4])+$signed(-{in[2003-:4],2'b0})+$signed(in[211-:4])+$signed(in[983-:4])+$signed(-in[1367-:4])+$signed(-{in[603-:4],2'b0})+$signed(-in[2011-:4])+$signed(-in[863-:4])+$signed(-in[227-:4])+$signed(-{in[1003-:4],2'b0})+$signed({in[363-:4],1'b0})+$signed(-in[1771-:4])+$signed(in[499-:4])+$signed(-in[375-:4])+$signed(-{in[639-:4],2'b0})+$signed(-{in[1279-:4],1'b0})+$signed(in[1663-:4])+$signed(sharing26)+$signed(-sharing27)+$signed(sharing38)+$signed(-sharing39)+$signed(sharing70)+$signed(-sharing71)+$signed(sharing108)+$signed(-sharing109)+$signed(sharing138)+$signed(sharing174)+$signed(-sharing175)+$signed(sharing199)+$signed(-sharing200)+$signed(-sharing206)+$signed(-sharing225)+$signed(0);
assign weighted_sum[16] = $signed({in[259-:4],1'b0})+$signed(-{in[1927-:4],1'b0})+$signed(-{in[523-:4],1'b0})+$signed(in[1167-:4])+$signed(in[1039-:4])+$signed(-in[667-:4])+$signed({in[927-:4],1'b0})+$signed(-in[163-:4])+$signed(in[1063-:4])+$signed({in[1195-:4],1'b0})+$signed(in[427-:4])+$signed(in[303-:4])+$signed(in[815-:4])+$signed(-in[435-:4])+$signed(in[1331-:4])+$signed(in[1843-:4])+$signed(-{in[951-:4],1'b0})+$signed(-{in[1987-:4],2'b0})+$signed({in[195-:4],1'b0})+$signed(in[67-:4])+$signed(-in[1347-:4])+$signed(-in[1475-:4])+$signed({in[1607-:4],1'b0})+$signed(in[1227-:4])+$signed(-{in[1619-:4],1'b0})+$signed({in[1495-:4],2'b0})+$signed(in[1371-:4])+$signed({in[95-:4],1'b0})+$signed(in[1887-:4])+$signed({in[1895-:4],1'b0})+$signed(-{in[2023-:4],1'b0})+$signed({in[879-:4],1'b0})+$signed(-in[243-:4])+$signed({in[1655-:4],2'b0})+$signed(in[1143-:4])+$signed({in[1659-:4],2'b0})+$signed({in[767-:4],1'b0})+$signed(sharing20)+$signed(sharing21)+$signed(sharing56)+$signed(-sharing57)+$signed(sharing80)+$signed(sharing81)+$signed(sharing112)+$signed(sharing113)+$signed(sharing139)+$signed(sharing140)+$signed(sharing164)+$signed(sharing191)+$signed(sharing209)+$signed(sharing221)+$signed(sharing222)+$signed(sharing244)+$signed(sharing253)+$signed(0);
assign weighted_sum[17] = $signed(-{in[1155-:4],1'b0})+$signed(in[899-:4])+$signed(in[891-:4])+$signed(-{in[1159-:4],2'b0})+$signed(-in[1671-:4])+$signed(-{in[1163-:4],3'b0})+$signed({in[1163-:4],1'b0})+$signed(-in[1419-:4])+$signed(-{in[1167-:4],3'b0})+$signed(-in[1807-:4])+$signed(-{in[1171-:4],3'b0})+$signed({in[1171-:4],1'b0})+$signed(-{in[1811-:4],1'b0})+$signed(-{in[1815-:4],2'b0})+$signed(-{in[1051-:4],2'b0})+$signed(-{in[931-:4],1'b0})+$signed(-in[1571-:4])+$signed(-{in[431-:4],3'b0})+$signed(-{in[1839-:4],3'b0})+$signed(in[1839-:4])+$signed(-{in[435-:4],3'b0})+$signed(-{in[1843-:4],3'b0})+$signed({in[435-:4],1'b0})+$signed(-{in[439-:4],2'b0})+$signed(in[439-:4])+$signed(-in[1975-:4])+$signed(-{in[1723-:4],2'b0})+$signed(in[187-:4])+$signed(in[63-:4])+$signed(in[191-:4])+$signed(-in[1343-:4])+$signed(in[1347-:4])+$signed(-in[1859-:4])+$signed(in[843-:4])+$signed(in[1739-:4])+$signed(-{in[1871-:4],2'b0})+$signed(-{in[1111-:4],2'b0})+$signed(in[1111-:4])+$signed(-{in[1759-:4],1'b0})+$signed(-in[1247-:4])+$signed(-{in[1763-:4],1'b0})+$signed(-{in[359-:4],2'b0})+$signed(-in[2023-:4])+$signed(-{in[491-:4],2'b0})+$signed(-{in[1003-:4],2'b0})+$signed(in[1771-:4])+$signed(in[367-:4])+$signed(-in[1007-:4])+$signed(-in[1775-:4])+$signed(-{in[371-:4],1'b0})+$signed(in[1267-:4])+$signed(-{in[375-:4],3'b0})+$signed(-{in[1779-:4],2'b0})+$signed(-{in[1783-:4],1'b0})+$signed(-{in[1915-:4],1'b0})+$signed(in[1659-:4])+$signed(in[1151-:4])+$signed(sharing22)+$signed(sharing23)+$signed(sharing50)+$signed(sharing51)+$signed(sharing82)+$signed(sharing83)+$signed(sharing114)+$signed(sharing115)+$signed(sharing141)+$signed(sharing142)+$signed(sharing165)+$signed(sharing194)+$signed(-sharing195)+$signed(sharing210)+$signed(sharing223)+$signed(sharing224)+$signed(sharing249)+$signed(0);
assign weighted_sum[18] = $signed(-{in[1923-:4],1'b0})+$signed(-in[1027-:4])+$signed(in[391-:4])+$signed({in[1291-:4],1'b0})+$signed(in[395-:4])+$signed(-{in[411-:4],1'b0})+$signed(-{in[795-:4],1'b0})+$signed(-in[1051-:4])+$signed(-in[35-:4])+$signed(-in[1187-:4])+$signed(-in[167-:4])+$signed(in[1579-:4])+$signed(in[1963-:4])+$signed(-{in[943-:4],1'b0})+$signed(in[1591-:4])+$signed(-in[1083-:4])+$signed(-{in[1087-:4],2'b0})+$signed(in[1215-:4])+$signed(-in[67-:4])+$signed(in[199-:4])+$signed(-in[711-:4])+$signed(-in[1351-:4])+$signed(-{in[1867-:4],1'b0})+$signed(-{in[1103-:4],2'b0})+$signed(in[1743-:4])+$signed({in[343-:4],1'b0})+$signed(in[859-:4])+$signed(in[347-:4])+$signed(in[611-:4])+$signed(in[231-:4])+$signed(-{in[1131-:4],1'b0})+$signed(-in[363-:4])+$signed(in[875-:4])+$signed(-{in[1135-:4],1'b0})+$signed(in[883-:4])+$signed(-in[503-:4])+$signed(sharing24)+$signed(sharing25)+$signed(sharing52)+$signed(sharing53)+$signed(sharing84)+$signed(sharing85)+$signed(sharing116)+$signed(sharing117)+$signed(sharing129)+$signed(-sharing130)+$signed(sharing166)+$signed(sharing167)+$signed(sharing183)+$signed(-sharing184)+$signed(sharing211)+$signed(sharing223)+$signed(-sharing224)+$signed(sharing233)+$signed(sharing244)+$signed(0);
assign weighted_sum[19] = $signed(-{in[643-:4],1'b0})+$signed(-in[515-:4])+$signed(in[1035-:4])+$signed(-{in[527-:4],1'b0})+$signed({in[1807-:4],1'b0})+$signed(-{in[1935-:4],1'b0})+$signed({in[1811-:4],1'b0})+$signed(-in[535-:4])+$signed(-{in[667-:4],2'b0})+$signed(in[1059-:4])+$signed(in[811-:4])+$signed(-{in[1583-:4],2'b0})+$signed(-{in[1587-:4],2'b0})+$signed(in[1075-:4])+$signed(-{in[567-:4],2'b0})+$signed(-in[1719-:4])+$signed(-{in[187-:4],1'b0})+$signed(-{in[1599-:4],2'b0})+$signed(-in[1343-:4])+$signed(in[1855-:4])+$signed(-{in[1987-:4],1'b0})+$signed(-in[195-:4])+$signed(in[451-:4])+$signed(-in[1995-:4])+$signed({in[847-:4],1'b0})+$signed(-in[591-:4])+$signed({in[1107-:4],1'b0})+$signed(-in[595-:4])+$signed(in[351-:4])+$signed(-{in[1639-:4],2'b0})+$signed(-in[363-:4])+$signed(in[1515-:4])+$signed(-in[1771-:4])+$signed({in[879-:4],1'b0})+$signed(in[1011-:4])+$signed(in[1139-:4])+$signed({in[1015-:4],1'b0})+$signed(-{in[1531-:4],2'b0})+$signed(sharing8)+$signed(-sharing9)+$signed(sharing54)+$signed(sharing55)+$signed(sharing86)+$signed(sharing87)+$signed(sharing118)+$signed(sharing119)+$signed(sharing143)+$signed(sharing144)+$signed(sharing168)+$signed(sharing187)+$signed(-sharing188)+$signed(sharing225)+$signed(sharing239)+$signed(-sharing241)+$signed(sharing250)+$signed(1);
assign weighted_sum[20] = $signed(-{in[1923-:4],1'b0})+$signed(in[1799-:4])+$signed({in[139-:4],1'b0})+$signed(-{in[1675-:4],1'b0})+$signed({in[1295-:4],1'b0})+$signed(-in[15-:4])+$signed(-in[399-:4])+$signed(-in[1679-:4])+$signed(-in[275-:4])+$signed(in[1427-:4])+$signed(-{in[1815-:4],1'b0})+$signed(in[895-:4])+$signed(-in[1823-:4])+$signed(-in[31-:4])+$signed(in[671-:4])+$signed({in[1699-:4],1'b0})+$signed(-in[163-:4])+$signed(in[935-:4])+$signed(-in[1195-:4])+$signed(-in[1971-:4])+$signed(-in[1207-:4])+$signed(-{in[571-:4],1'b0})+$signed(-in[827-:4])+$signed(-{in[1087-:4],1'b0})+$signed(in[967-:4])+$signed(in[1991-:4])+$signed(-in[1103-:4])+$signed({in[1495-:4],1'b0})+$signed(in[87-:4])+$signed({in[1243-:4],1'b0})+$signed(-in[1131-:4])+$signed(-{in[495-:4],1'b0})+$signed(-in[1135-:4])+$signed(in[1647-:4])+$signed(in[1271-:4])+$signed({in[1659-:4],1'b0})+$signed(-in[635-:4])+$signed(in[1535-:4])+$signed(sharing22)+$signed(-sharing23)+$signed(sharing34)+$signed(-sharing35)+$signed(sharing90)+$signed(-sharing91)+$signed(sharing122)+$signed(-sharing123)+$signed(sharing145)+$signed(sharing146)+$signed(sharing169)+$signed(sharing192)+$signed(-sharing211)+$signed(-sharing219)+$signed(sharing237)+$signed(sharing240)+$signed(-2);
assign weighted_sum[21] = $signed(-in[891-:4])+$signed(in[1931-:4])+$signed(-{in[1679-:4],1'b0})+$signed(-{in[1807-:4],1'b0})+$signed(-in[399-:4])+$signed(-{in[767-:4],1'b0})+$signed({in[1427-:4],1'b0})+$signed(-{in[1567-:4],2'b0})+$signed(-{in[1823-:4],1'b0})+$signed(-in[1695-:4])+$signed(in[1059-:4])+$signed(-{in[1707-:4],2'b0})+$signed({in[1971-:4],2'b0})+$signed(-in[1203-:4])+$signed(in[1079-:4])+$signed(in[183-:4])+$signed({in[1339-:4],1'b0})+$signed(in[827-:4])+$signed(in[1595-:4])+$signed({in[1343-:4],1'b0})+$signed(-in[451-:4])+$signed({in[1863-:4],1'b0})+$signed(-in[455-:4])+$signed(in[1103-:4])+$signed(in[1487-:4])+$signed(-in[1623-:4])+$signed(-{in[1755-:4],2'b0})+$signed(-{in[1627-:4],1'b0})+$signed({in[1247-:4],1'b0})+$signed(-{in[1759-:4],1'b0})+$signed({in[611-:4],1'b0})+$signed(-{in[1771-:4],1'b0})+$signed(-{in[751-:4],1'b0})+$signed(-in[111-:4])+$signed(-in[251-:4])+$signed(in[1903-:4])+$signed({in[1907-:4],1'b0})+$signed(-in[1651-:4])+$signed(in[1015-:4])+$signed({in[1915-:4],2'b0})+$signed(in[1787-:4])+$signed({in[1919-:4],2'b0})+$signed({in[383-:4],1'b0})+$signed(sharing26)+$signed(sharing27)+$signed(sharing62)+$signed(-sharing63)+$signed(sharing88)+$signed(-sharing89)+$signed(sharing110)+$signed(-sharing111)+$signed(sharing136)+$signed(-sharing137)+$signed(sharing156)+$signed(-sharing157)+$signed(sharing181)+$signed(-sharing182)+$signed(sharing201)+$signed(sharing229)+$signed(sharing246)+$signed(2);
assign weighted_sum[22] = $signed({in[1539-:4],1'b0})+$signed(in[515-:4])+$signed({in[903-:4],1'b0})+$signed(-in[7-:4])+$signed({in[907-:4],1'b0})+$signed({in[911-:4],2'b0})+$signed(in[1807-:4])+$signed({in[403-:4],1'b0})+$signed(in[915-:4])+$signed({in[411-:4],1'b0})+$signed(in[1051-:4])+$signed(-in[163-:4])+$signed(-in[295-:4])+$signed(in[1963-:4])+$signed({in[179-:4],1'b0})+$signed(-in[51-:4])+$signed(in[563-:4])+$signed({in[1591-:4],1'b0})+$signed({in[1083-:4],1'b0})+$signed({in[1851-:4],1'b0})+$signed({in[1855-:4],1'b0})+$signed(-in[319-:4])+$signed(in[1087-:4])+$signed(in[451-:4])+$signed({in[455-:4],1'b0})+$signed({in[855-:4],2'b0})+$signed({in[1879-:4],1'b0})+$signed({in[859-:4],2'b0})+$signed(in[1499-:4])+$signed({in[351-:4],1'b0})+$signed({in[355-:4],1'b0})+$signed({in[231-:4],1'b0})+$signed(-in[1639-:4])+$signed(in[1767-:4])+$signed(in[1895-:4])+$signed(-in[111-:4])+$signed({in[1139-:4],1'b0})+$signed(in[499-:4])+$signed(in[1911-:4])+$signed({in[511-:4],1'b0})+$signed(sharing10)+$signed(-sharing11)+$signed(sharing46)+$signed(-sharing47)+$signed(sharing74)+$signed(-sharing75)+$signed(sharing96)+$signed(-sharing97)+$signed(sharing132)+$signed(-sharing133)+$signed(sharing170)+$signed(sharing171)+$signed(sharing193)+$signed(sharing207)+$signed(-sharing208)+$signed(0);
assign weighted_sum[23] = $signed({in[1027-:4],2'b0})+$signed({in[1031-:4],2'b0})+$signed(-in[1415-:4])+$signed(-in[775-:4])+$signed(in[135-:4])+$signed(in[651-:4])+$signed(in[1675-:4])+$signed(-in[1551-:4])+$signed(-{in[1555-:4],1'b0})+$signed({in[1567-:4],1'b0})+$signed(-in[31-:4])+$signed({in[799-:4],1'b0})+$signed(-in[671-:4])+$signed({in[1571-:4],1'b0})+$signed(-in[1187-:4])+$signed(-{in[39-:4],1'b0})+$signed({in[295-:4],1'b0})+$signed({in[299-:4],2'b0})+$signed(-in[1451-:4])+$signed(in[1579-:4])+$signed(in[1203-:4])+$signed(-in[823-:4])+$signed({in[955-:4],1'b0})+$signed({in[1471-:4],1'b0})+$signed(-in[63-:4])+$signed(-in[1599-:4])+$signed(-in[203-:4])+$signed(in[1483-:4])+$signed({in[975-:4],2'b0})+$signed(-{in[207-:4],1'b0})+$signed({in[851-:4],2'b0})+$signed(in[471-:4])+$signed(-{in[95-:4],2'b0})+$signed(in[1759-:4])+$signed(-in[99-:4])+$signed(-in[239-:4])+$signed(-in[755-:4])+$signed(-in[503-:4])+$signed(in[1019-:4])+$signed({in[1023-:4],2'b0})+$signed({in[639-:4],1'b0})+$signed(in[511-:4])+$signed(sharing16)+$signed(-sharing17)+$signed(sharing42)+$signed(-sharing43)+$signed(sharing64)+$signed(-sharing65)+$signed(sharing118)+$signed(-sharing119)+$signed(sharing131)+$signed(sharing176)+$signed(-sharing193)+$signed(-sharing251)+$signed(-sharing253)+$signed(1);
assign weighted_sum[24] = $signed(-{in[1159-:4],1'b0})+$signed(-{in[1031-:4],1'b0})+$signed(-in[523-:4])+$signed(in[779-:4])+$signed({in[527-:4],1'b0})+$signed(in[1935-:4])+$signed(in[1687-:4])+$signed(in[803-:4])+$signed(in[1443-:4])+$signed(in[1447-:4])+$signed({in[1075-:4],1'b0})+$signed(-{in[1079-:4],1'b0})+$signed(in[951-:4])+$signed(-{in[1083-:4],1'b0})+$signed({in[1987-:4],1'b0})+$signed(-in[207-:4])+$signed(in[847-:4])+$signed(in[83-:4])+$signed(in[1875-:4])+$signed(-{in[983-:4],2'b0})+$signed(in[1751-:4])+$signed(in[1627-:4])+$signed(in[1503-:4])+$signed(-in[227-:4])+$signed(-{in[1767-:4],1'b0})+$signed(in[1639-:4])+$signed(-{in[619-:4],2'b0})+$signed(-in[1003-:4])+$signed(in[1259-:4])+$signed(in[1387-:4])+$signed(in[1907-:4])+$signed(-in[383-:4])+$signed(sharing28)+$signed(sharing29)+$signed(sharing56)+$signed(sharing57)+$signed(sharing88)+$signed(sharing89)+$signed(sharing120)+$signed(sharing121)+$signed(sharing147)+$signed(sharing148)+$signed(sharing172)+$signed(sharing194)+$signed(sharing195)+$signed(sharing212)+$signed(sharing213)+$signed(sharing226)+$signed(sharing234)+$signed(sharing239)+$signed(sharing245)+$signed(sharing251)+$signed(2);
assign weighted_sum[25] = $signed({in[1019-:4],1'b0})+$signed(-in[3-:4])+$signed({in[139-:4],2'b0})+$signed({in[1935-:4],1'b0})+$signed(-in[1687-:4])+$signed(-in[663-:4])+$signed(-in[1319-:4])+$signed(in[1703-:4])+$signed(-in[299-:4])+$signed({in[1839-:4],2'b0})+$signed({in[1967-:4],1'b0})+$signed({in[1843-:4],2'b0})+$signed({in[567-:4],1'b0})+$signed(-{in[1723-:4],1'b0})+$signed(in[1851-:4])+$signed({in[1855-:4],1'b0})+$signed({in[1859-:4],1'b0})+$signed({in[583-:4],1'b0})+$signed(in[199-:4])+$signed(in[1995-:4])+$signed(in[1883-:4])+$signed({in[1891-:4],2'b0})+$signed(-in[1123-:4])+$signed({in[1895-:4],2'b0})+$signed(in[1767-:4])+$signed(-{in[1267-:4],1'b0})+$signed(in[755-:4])+$signed({in[1911-:4],1'b0})+$signed({in[507-:4],1'b0})+$signed({in[1663-:4],1'b0})+$signed(-in[639-:4])+$signed(sharing2)+$signed(-sharing3)+$signed(sharing58)+$signed(sharing59)+$signed(sharing90)+$signed(sharing91)+$signed(sharing112)+$signed(-sharing113)+$signed(sharing141)+$signed(-sharing142)+$signed(sharing172)+$signed(sharing196)+$signed(sharing197)+$signed(sharing227)+$signed(sharing246)+$signed(sharing252)+$signed(sharing254)+$signed(sharing255)+$signed(0);
assign weighted_sum[26] = $signed(-in[387-:4])+$signed(-{in[1031-:4],1'b0})+$signed(in[383-:4])+$signed(-{in[1171-:4],1'b0})+$signed(in[1555-:4])+$signed({in[919-:4],1'b0})+$signed(-{in[927-:4],1'b0})+$signed({in[671-:4],1'b0})+$signed(in[1279-:4])+$signed({in[1447-:4],1'b0})+$signed(in[43-:4])+$signed(in[431-:4])+$signed(in[815-:4])+$signed(in[307-:4])+$signed(in[955-:4])+$signed(-in[1855-:4])+$signed(-in[971-:4])+$signed(-{in[975-:4],1'b0})+$signed(-{in[979-:4],1'b0})+$signed(in[2003-:4])+$signed(-in[343-:4])+$signed(-{in[1627-:4],1'b0})+$signed({in[1503-:4],1'b0})+$signed(-in[1759-:4])+$signed(-{in[1767-:4],2'b0})+$signed(-in[1383-:4])+$signed(-in[2027-:4])+$signed({in[755-:4],1'b0})+$signed({in[1011-:4],1'b0})+$signed({in[1651-:4],1'b0})+$signed({in[1015-:4],2'b0})+$signed({in[759-:4],1'b0})+$signed(in[375-:4])+$signed({in[1779-:4],1'b0})+$signed({in[635-:4],1'b0})+$signed({in[1787-:4],1'b0})+$signed(-{in[1023-:4],1'b0})+$signed(in[1791-:4])+$signed(sharing6)+$signed(-sharing7)+$signed(sharing58)+$signed(-sharing59)+$signed(sharing66)+$signed(-sharing67)+$signed(sharing122)+$signed(sharing123)+$signed(sharing149)+$signed(sharing150)+$signed(sharing166)+$signed(-sharing167)+$signed(sharing198)+$signed(sharing214)+$signed(sharing215)+$signed(sharing228)+$signed(sharing235)+$signed(3);
assign weighted_sum[27] = $signed({in[1795-:4],2'b0})+$signed({in[1155-:4],1'b0})+$signed(in[771-:4])+$signed({in[395-:4],1'b0})+$signed(in[399-:4])+$signed({in[1555-:4],1'b0})+$signed(in[1559-:4])+$signed(-in[1047-:4])+$signed({in[155-:4],1'b0})+$signed(-{in[411-:4],1'b0})+$signed(-in[283-:4])+$signed(-in[543-:4])+$signed(in[1067-:4])+$signed(in[1963-:4])+$signed(in[559-:4])+$signed(in[1583-:4])+$signed({in[1975-:4],1'b0})+$signed({in[1851-:4],1'b0})+$signed({in[831-:4],1'b0})+$signed({in[447-:4],1'b0})+$signed(-in[1983-:4])+$signed(-in[579-:4])+$signed(-in[963-:4])+$signed(in[1603-:4])+$signed(-{in[843-:4],1'b0})+$signed(-in[1099-:4])+$signed({in[1747-:4],1'b0})+$signed(in[855-:4])+$signed(-in[1623-:4])+$signed(-in[603-:4])+$signed(-in[1883-:4])+$signed({in[1119-:4],1'b0})+$signed({in[2015-:4],1'b0})+$signed({in[2019-:4],1'b0})+$signed(in[615-:4])+$signed({in[619-:4],1'b0})+$signed({in[1259-:4],1'b0})+$signed(-in[1643-:4])+$signed(-{in[1771-:4],1'b0})+$signed(-in[1011-:4])+$signed(-in[1139-:4])+$signed({in[1919-:4],1'b0})+$signed(in[1663-:4])+$signed(sharing28)+$signed(-sharing29)+$signed(sharing60)+$signed(sharing61)+$signed(sharing80)+$signed(-sharing81)+$signed(sharing124)+$signed(sharing125)+$signed(sharing173)+$signed(sharing216)+$signed(sharing247)+$signed(0);
assign weighted_sum[28] = $signed(-{in[259-:4],2'b0})+$signed(in[1031-:4])+$signed(-in[903-:4])+$signed(in[651-:4])+$signed(in[1419-:4])+$signed(in[1295-:4])+$signed(in[1679-:4])+$signed(in[1935-:4])+$signed({in[915-:4],1'b0})+$signed(in[1299-:4])+$signed(-{in[1559-:4],2'b0})+$signed(in[795-:4])+$signed({in[187-:4],2'b0})+$signed({in[191-:4],1'b0})+$signed(-in[959-:4])+$signed(-in[1215-:4])+$signed(in[323-:4])+$signed(-{in[1611-:4],2'b0})+$signed(in[1867-:4])+$signed(-{in[207-:4],2'b0})+$signed({in[1871-:4],1'b0})+$signed(-in[975-:4])+$signed(in[1619-:4])+$signed(in[1623-:4])+$signed(-in[1755-:4])+$signed(-in[95-:4])+$signed({in[867-:4],1'b0})+$signed(in[867-:4])+$signed({in[1635-:4],1'b0})+$signed({in[1639-:4],1'b0})+$signed(in[1895-:4])+$signed(-{in[1519-:4],1'b0})+$signed(-{in[1523-:4],1'b0})+$signed(-in[1655-:4])+$signed({in[1019-:4],1'b0})+$signed(-in[1659-:4])+$signed(sharing20)+$signed(-sharing21)+$signed(sharing40)+$signed(-sharing41)+$signed(sharing92)+$signed(sharing93)+$signed(sharing126)+$signed(sharing149)+$signed(-sharing150)+$signed(-sharing168)+$signed(sharing199)+$signed(sharing200)+$signed(sharing202)+$signed(sharing229)+$signed(sharing242)+$signed(1);
assign weighted_sum[29] = $signed(-in[1539-:4])+$signed(in[771-:4])+$signed(in[1667-:4])+$signed(in[1803-:4])+$signed(in[1163-:4])+$signed(-{in[527-:4],2'b0})+$signed({in[271-:4],1'b0})+$signed(in[527-:4])+$signed({in[1679-:4],2'b0})+$signed(in[1679-:4])+$signed({in[1555-:4],1'b0})+$signed({in[1683-:4],2'b0})+$signed({in[279-:4],2'b0})+$signed({in[1559-:4],1'b0})+$signed({in[283-:4],3'b0})+$signed(in[1951-:4])+$signed(-in[299-:4])+$signed(in[1195-:4])+$signed(-in[1967-:4])+$signed(-{in[1591-:4],1'b0})+$signed(-in[1207-:4])+$signed(in[1463-:4])+$signed({in[1723-:4],1'b0})+$signed({in[963-:4],2'b0})+$signed(-in[1475-:4])+$signed({in[327-:4],2'b0})+$signed({in[967-:4],1'b0})+$signed(in[967-:4])+$signed(-in[587-:4])+$signed(-{in[79-:4],1'b0})+$signed(-{in[1875-:4],1'b0})+$signed(-{in[87-:4],1'b0})+$signed(-in[855-:4])+$signed(-in[475-:4])+$signed(-in[219-:4])+$signed(in[995-:4])+$signed({in[1639-:4],2'b0})+$signed(-{in[2027-:4],1'b0})+$signed({in[1007-:4],2'b0})+$signed(-in[879-:4])+$signed(in[1139-:4])+$signed(sharing14)+$signed(-sharing15)+$signed(sharing62)+$signed(sharing63)+$signed(sharing68)+$signed(-sharing69)+$signed(sharing120)+$signed(-sharing121)+$signed(sharing151)+$signed(sharing152)+$signed(sharing174)+$signed(sharing175)+$signed(-sharing203)+$signed(sharing228)+$signed(-sharing230)+$signed(2);
assign weighted_sum[30] = $signed(-in[515-:4])+$signed(-{in[775-:4],1'b0})+$signed(-in[519-:4])+$signed({in[1035-:4],1'b0})+$signed(-in[651-:4])+$signed(-in[1291-:4])+$signed(-{in[1551-:4],2'b0})+$signed(-{in[151-:4],1'b0})+$signed(-{in[1687-:4],1'b0})+$signed({in[1051-:4],1'b0})+$signed(-in[283-:4])+$signed({in[1311-:4],1'b0})+$signed({in[1315-:4],1'b0})+$signed(-{in[935-:4],1'b0})+$signed(-{in[1703-:4],1'b0})+$signed({in[947-:4],1'b0})+$signed(-in[819-:4])+$signed(-{in[1715-:4],1'b0})+$signed({in[951-:4],1'b0})+$signed(-{in[1975-:4],1'b0})+$signed(-in[1339-:4])+$signed(-in[1595-:4])+$signed(-{in[1599-:4],1'b0})+$signed(-{in[1603-:4],2'b0})+$signed(-{in[1219-:4],1'b0})+$signed(-{in[1607-:4],2'b0})+$signed(-in[331-:4])+$signed(-{in[207-:4],1'b0})+$signed({in[215-:4],1'b0})+$signed({in[1623-:4],1'b0})+$signed(-{in[987-:4],2'b0})+$signed(in[219-:4])+$signed(-in[2011-:4])+$signed(-{in[99-:4],2'b0})+$signed(-{in[867-:4],1'b0})+$signed(-{in[1123-:4],1'b0})+$signed(in[1767-:4])+$signed(-in[619-:4])+$signed({in[1007-:4],1'b0})+$signed(in[111-:4])+$signed(-in[1903-:4])+$signed(-{in[883-:4],1'b0})+$signed(in[243-:4])+$signed(-{in[1659-:4],2'b0})+$signed(-{in[1663-:4],2'b0})+$signed(in[1535-:4])+$signed(sharing30)+$signed(sharing31)+$signed(sharing52)+$signed(-sharing53)+$signed(sharing94)+$signed(sharing95)+$signed(sharing114)+$signed(-sharing115)+$signed(sharing153)+$signed(sharing154)+$signed(-sharing169)+$signed(sharing178)+$signed(-sharing179)+$signed(sharing214)+$signed(-sharing215)+$signed(-sharing227)+$signed(1);
assign weighted_sum[31] = $signed(-in[1035-:4])+$signed(-in[1675-:4])+$signed({in[1935-:4],1'b0})+$signed(-{in[1551-:4],1'b0})+$signed(-in[143-:4])+$signed(in[1555-:4])+$signed({in[919-:4],1'b0})+$signed({in[1175-:4],1'b0})+$signed({in[923-:4],2'b0})+$signed(-in[155-:4])+$signed({in[927-:4],2'b0})+$signed({in[931-:4],1'b0})+$signed(in[1827-:4])+$signed(in[1323-:4])+$signed(-in[303-:4])+$signed(-{in[307-:4],1'b0})+$signed(in[951-:4])+$signed(in[1335-:4])+$signed(-in[1975-:4])+$signed({in[447-:4],1'b0})+$signed(-in[703-:4])+$signed({in[579-:4],1'b0})+$signed(in[195-:4])+$signed({in[1475-:4],1'b0})+$signed({in[967-:4],2'b0})+$signed(in[979-:4])+$signed(in[1879-:4])+$signed(-in[223-:4])+$signed(in[1887-:4])+$signed(-{in[99-:4],1'b0})+$signed(-in[355-:4])+$signed({in[1127-:4],1'b0})+$signed(-in[359-:4])+$signed({in[239-:4],1'b0})+$signed(in[239-:4])+$signed(in[495-:4])+$signed({in[243-:4],2'b0})+$signed({in[115-:4],1'b0})+$signed(-in[623-:4])+$signed(-{in[1655-:4],1'b0})+$signed(in[1271-:4])+$signed({in[251-:4],1'b0})+$signed(in[1275-:4])+$signed({in[255-:4],1'b0})+$signed(sharing30)+$signed(-sharing31)+$signed(sharing44)+$signed(-sharing45)+$signed(sharing84)+$signed(-sharing85)+$signed(sharing102)+$signed(-sharing103)+$signed(sharing151)+$signed(-sharing152)+$signed(sharing176)+$signed(-sharing198)+$signed(2);
assign relu_out[0] = (weighted_sum[0][9]==1) ? 4'd0 : (weighted_sum[0][8:2] > 6 ? 4'd6 : weighted_sum[0][5:2]);
assign relu_out[1] = (weighted_sum[1][9]==1) ? 4'd0 : (weighted_sum[1][8:2] > 6 ? 4'd6 : weighted_sum[1][5:2]);
assign relu_out[2] = (weighted_sum[2][9]==1) ? 4'd0 : (weighted_sum[2][8:2] > 6 ? 4'd6 : weighted_sum[2][5:2]);
assign relu_out[3] = (weighted_sum[3][9]==1) ? 4'd0 : (weighted_sum[3][8:2] > 6 ? 4'd6 : weighted_sum[3][5:2]);
assign relu_out[4] = (weighted_sum[4][9]==1) ? 4'd0 : (weighted_sum[4][8:2] > 6 ? 4'd6 : weighted_sum[4][5:2]);
assign relu_out[5] = (weighted_sum[5][9]==1) ? 4'd0 : (weighted_sum[5][8:2] > 6 ? 4'd6 : weighted_sum[5][5:2]);
assign relu_out[6] = (weighted_sum[6][9]==1) ? 4'd0 : (weighted_sum[6][8:2] > 6 ? 4'd6 : weighted_sum[6][5:2]);
assign relu_out[7] = (weighted_sum[7][9]==1) ? 4'd0 : (weighted_sum[7][8:2] > 6 ? 4'd6 : weighted_sum[7][5:2]);
assign relu_out[8] = (weighted_sum[8][9]==1) ? 4'd0 : (weighted_sum[8][8:2] > 6 ? 4'd6 : weighted_sum[8][5:2]);
assign relu_out[9] = (weighted_sum[9][9]==1) ? 4'd0 : (weighted_sum[9][8:2] > 6 ? 4'd6 : weighted_sum[9][5:2]);
assign relu_out[10] = (weighted_sum[10][9]==1) ? 4'd0 : (weighted_sum[10][8:2] > 6 ? 4'd6 : weighted_sum[10][5:2]);
assign relu_out[11] = (weighted_sum[11][9]==1) ? 4'd0 : (weighted_sum[11][8:2] > 6 ? 4'd6 : weighted_sum[11][5:2]);
assign relu_out[12] = (weighted_sum[12][9]==1) ? 4'd0 : (weighted_sum[12][8:2] > 6 ? 4'd6 : weighted_sum[12][5:2]);
assign relu_out[13] = (weighted_sum[13][9]==1) ? 4'd0 : (weighted_sum[13][8:2] > 6 ? 4'd6 : weighted_sum[13][5:2]);
assign relu_out[14] = (weighted_sum[14][9]==1) ? 4'd0 : (weighted_sum[14][8:2] > 6 ? 4'd6 : weighted_sum[14][5:2]);
assign relu_out[15] = (weighted_sum[15][9]==1) ? 4'd0 : (weighted_sum[15][8:2] > 6 ? 4'd6 : weighted_sum[15][5:2]);
assign relu_out[16] = (weighted_sum[16][9]==1) ? 4'd0 : (weighted_sum[16][8:2] > 6 ? 4'd6 : weighted_sum[16][5:2]);
assign relu_out[17] = (weighted_sum[17][9]==1) ? 4'd0 : (weighted_sum[17][8:2] > 6 ? 4'd6 : weighted_sum[17][5:2]);
assign relu_out[18] = (weighted_sum[18][9]==1) ? 4'd0 : (weighted_sum[18][8:2] > 6 ? 4'd6 : weighted_sum[18][5:2]);
assign relu_out[19] = (weighted_sum[19][9]==1) ? 4'd0 : (weighted_sum[19][8:2] > 6 ? 4'd6 : weighted_sum[19][5:2]);
assign relu_out[20] = (weighted_sum[20][9]==1) ? 4'd0 : (weighted_sum[20][8:2] > 6 ? 4'd6 : weighted_sum[20][5:2]);
assign relu_out[21] = (weighted_sum[21][9]==1) ? 4'd0 : (weighted_sum[21][8:2] > 6 ? 4'd6 : weighted_sum[21][5:2]);
assign relu_out[22] = (weighted_sum[22][9]==1) ? 4'd0 : (weighted_sum[22][8:2] > 6 ? 4'd6 : weighted_sum[22][5:2]);
assign relu_out[23] = (weighted_sum[23][9]==1) ? 4'd0 : (weighted_sum[23][8:2] > 6 ? 4'd6 : weighted_sum[23][5:2]);
assign relu_out[24] = (weighted_sum[24][9]==1) ? 4'd0 : (weighted_sum[24][8:2] > 6 ? 4'd6 : weighted_sum[24][5:2]);
assign relu_out[25] = (weighted_sum[25][9]==1) ? 4'd0 : (weighted_sum[25][8:2] > 6 ? 4'd6 : weighted_sum[25][5:2]);
assign relu_out[26] = (weighted_sum[26][9]==1) ? 4'd0 : (weighted_sum[26][8:2] > 6 ? 4'd6 : weighted_sum[26][5:2]);
assign relu_out[27] = (weighted_sum[27][9]==1) ? 4'd0 : (weighted_sum[27][8:2] > 6 ? 4'd6 : weighted_sum[27][5:2]);
assign relu_out[28] = (weighted_sum[28][9]==1) ? 4'd0 : (weighted_sum[28][8:2] > 6 ? 4'd6 : weighted_sum[28][5:2]);
assign relu_out[29] = (weighted_sum[29][9]==1) ? 4'd0 : (weighted_sum[29][8:2] > 6 ? 4'd6 : weighted_sum[29][5:2]);
assign relu_out[30] = (weighted_sum[30][9]==1) ? 4'd0 : (weighted_sum[30][8:2] > 6 ? 4'd6 : weighted_sum[30][5:2]);
assign relu_out[31] = (weighted_sum[31][9]==1) ? 4'd0 : (weighted_sum[31][8:2] > 6 ? 4'd6 : weighted_sum[31][5:2]);
assign out = {relu_out[31],relu_out[30],relu_out[29],relu_out[28],relu_out[27],relu_out[26],relu_out[25],relu_out[24],relu_out[23],relu_out[22],relu_out[21],relu_out[20],relu_out[19],relu_out[18],relu_out[17],relu_out[16],relu_out[15],relu_out[14],relu_out[13],relu_out[12],relu_out[11],relu_out[10],relu_out[9],relu_out[8],relu_out[7],relu_out[6],relu_out[5],relu_out[4],relu_out[3],relu_out[2],relu_out[1],relu_out[0]};

endmodule
