module conv1 (
	input [6271:0] in,
	output [2027:0] out
);

wire [3:0] relu_out [0:506];
wire [12:0] weighted_sum [0:506];
wire [12:0] sharing0;
wire [12:0] sharing1;
wire [12:0] sharing2;
wire [12:0] sharing3;
wire [12:0] sharing4;
wire [12:0] sharing5;
wire [12:0] sharing6;
wire [12:0] sharing7;
wire [12:0] sharing8;
wire [12:0] sharing9;
wire [12:0] sharing10;
wire [12:0] sharing11;
wire [12:0] sharing12;
wire [12:0] sharing13;
wire [12:0] sharing14;
wire [12:0] sharing15;
wire [12:0] sharing16;
wire [12:0] sharing17;
wire [12:0] sharing18;
wire [12:0] sharing19;
wire [12:0] sharing20;
wire [12:0] sharing21;
wire [12:0] sharing22;
wire [12:0] sharing23;
wire [12:0] sharing24;
wire [12:0] sharing25;
wire [12:0] sharing26;
wire [12:0] sharing27;
wire [12:0] sharing28;
wire [12:0] sharing29;
wire [12:0] sharing30;
wire [12:0] sharing31;
wire [12:0] sharing32;
wire [12:0] sharing33;
wire [12:0] sharing34;
wire [12:0] sharing35;
wire [12:0] sharing36;
wire [12:0] sharing37;
wire [12:0] sharing38;
wire [12:0] sharing39;
wire [12:0] sharing40;
wire [12:0] sharing41;
wire [12:0] sharing42;
wire [12:0] sharing43;
wire [12:0] sharing44;
wire [12:0] sharing45;
wire [12:0] sharing46;
wire [12:0] sharing47;
wire [12:0] sharing48;
wire [12:0] sharing49;
wire [12:0] sharing50;
wire [12:0] sharing51;
wire [12:0] sharing52;
wire [12:0] sharing53;
wire [12:0] sharing54;
wire [12:0] sharing55;
wire [12:0] sharing56;
wire [12:0] sharing57;
wire [12:0] sharing58;
wire [12:0] sharing59;
wire [12:0] sharing60;
wire [12:0] sharing61;
wire [12:0] sharing62;
wire [12:0] sharing63;
wire [12:0] sharing64;
wire [12:0] sharing65;
wire [12:0] sharing66;
wire [12:0] sharing67;
wire [12:0] sharing68;
wire [12:0] sharing69;
wire [12:0] sharing70;
wire [12:0] sharing71;
wire [12:0] sharing72;
wire [12:0] sharing73;
wire [12:0] sharing74;
wire [12:0] sharing75;
wire [12:0] sharing76;
wire [12:0] sharing77;
wire [12:0] sharing78;
wire [12:0] sharing79;
wire [12:0] sharing80;
wire [12:0] sharing81;
wire [12:0] sharing82;
wire [12:0] sharing83;
wire [12:0] sharing84;
wire [12:0] sharing85;
wire [12:0] sharing86;
wire [12:0] sharing87;
wire [12:0] sharing88;
wire [12:0] sharing89;
wire [12:0] sharing90;
wire [12:0] sharing91;
wire [12:0] sharing92;
wire [12:0] sharing93;
wire [12:0] sharing94;
wire [12:0] sharing95;
wire [12:0] sharing96;
wire [12:0] sharing97;
wire [12:0] sharing98;
wire [12:0] sharing99;
wire [12:0] sharing100;
wire [12:0] sharing101;
wire [12:0] sharing102;
wire [12:0] sharing103;
wire [12:0] sharing104;
wire [12:0] sharing105;
wire [12:0] sharing106;
wire [12:0] sharing107;
wire [12:0] sharing108;
wire [12:0] sharing109;
wire [12:0] sharing110;
wire [12:0] sharing111;
wire [12:0] sharing112;
wire [12:0] sharing113;
wire [12:0] sharing114;
wire [12:0] sharing115;
wire [12:0] sharing116;
wire [12:0] sharing117;
wire [12:0] sharing118;
wire [12:0] sharing119;
wire [12:0] sharing120;
wire [12:0] sharing121;
wire [12:0] sharing122;
wire [12:0] sharing123;
wire [12:0] sharing124;
wire [12:0] sharing125;
wire [12:0] sharing126;
wire [12:0] sharing127;
wire [12:0] sharing128;
wire [12:0] sharing129;
wire [12:0] sharing130;
wire [12:0] sharing131;
wire [12:0] sharing132;
wire [12:0] sharing133;
wire [12:0] sharing134;
wire [12:0] sharing135;
wire [12:0] sharing136;
wire [12:0] sharing137;
wire [12:0] sharing138;
wire [12:0] sharing139;
wire [12:0] sharing140;
wire [12:0] sharing141;
wire [12:0] sharing142;
wire [12:0] sharing143;
wire [12:0] sharing144;
wire [12:0] sharing145;
wire [12:0] sharing146;
wire [12:0] sharing147;
wire [12:0] sharing148;
wire [12:0] sharing149;
wire [12:0] sharing150;
wire [12:0] sharing151;
wire [12:0] sharing152;
wire [12:0] sharing153;
wire [12:0] sharing154;
wire [12:0] sharing155;
wire [12:0] sharing156;
wire [12:0] sharing157;
wire [12:0] sharing158;
wire [12:0] sharing159;
wire [12:0] sharing160;
wire [12:0] sharing161;
wire [12:0] sharing162;
wire [12:0] sharing163;
wire [12:0] sharing164;
wire [12:0] sharing165;
wire [12:0] sharing166;
wire [12:0] sharing167;
wire [12:0] sharing168;

assign sharing0 = $signed({in[7-:8],2'b0})+$signed(in[7-:8])+$signed({in[15-:8],2'b0})+$signed(in[463-:8]);
assign sharing1 = $signed({in[23-:8],2'b0})+$signed(in[23-:8])+$signed({in[31-:8],2'b0})+$signed(in[479-:8]);
assign sharing2 = $signed({in[39-:8],2'b0})+$signed(in[39-:8])+$signed({in[47-:8],2'b0})+$signed(in[495-:8]);
assign sharing3 = $signed({in[55-:8],2'b0})+$signed(in[55-:8])+$signed({in[63-:8],2'b0})+$signed(in[511-:8]);
assign sharing4 = $signed({in[71-:8],2'b0})+$signed(in[71-:8])+$signed({in[79-:8],2'b0})+$signed(in[527-:8]);
assign sharing5 = $signed({in[87-:8],2'b0})+$signed(in[87-:8])+$signed({in[95-:8],2'b0})+$signed(in[543-:8]);
assign sharing6 = $signed({in[119-:8],2'b0})+$signed(in[119-:8])+$signed({in[127-:8],2'b0})+$signed(in[575-:8]);
assign sharing7 = $signed({in[135-:8],2'b0})+$signed(in[135-:8])+$signed({in[143-:8],2'b0})+$signed(in[591-:8]);
assign sharing8 = $signed({in[151-:8],2'b0})+$signed(in[151-:8])+$signed({in[159-:8],2'b0})+$signed(in[607-:8]);
assign sharing9 = $signed({in[167-:8],2'b0})+$signed(in[167-:8])+$signed({in[175-:8],2'b0})+$signed(in[623-:8]);
assign sharing10 = $signed({in[183-:8],2'b0})+$signed(in[183-:8])+$signed({in[191-:8],2'b0})+$signed(in[639-:8]);
assign sharing11 = $signed({in[199-:8],2'b0})+$signed(in[199-:8])+$signed({in[207-:8],2'b0})+$signed(in[655-:8]);
assign sharing12 = $signed({in[455-:8],2'b0})+$signed(in[455-:8])+$signed({in[463-:8],2'b0})+$signed(in[911-:8]);
assign sharing13 = $signed({in[487-:8],2'b0})+$signed(in[487-:8])+$signed({in[495-:8],2'b0})+$signed(in[943-:8]);
assign sharing14 = $signed({in[503-:8],2'b0})+$signed(in[503-:8])+$signed({in[511-:8],2'b0})+$signed(in[959-:8]);
assign sharing15 = $signed({in[519-:8],2'b0})+$signed(in[519-:8])+$signed({in[527-:8],2'b0})+$signed(in[975-:8]);
assign sharing16 = $signed({in[535-:8],2'b0})+$signed(in[535-:8])+$signed({in[543-:8],2'b0})+$signed(in[991-:8]);
assign sharing17 = $signed({in[551-:8],2'b0})+$signed(in[551-:8])+$signed({in[559-:8],2'b0})+$signed(in[1007-:8]);
assign sharing18 = $signed({in[567-:8],2'b0})+$signed(in[567-:8])+$signed({in[575-:8],2'b0})+$signed(in[1023-:8]);
assign sharing19 = $signed({in[583-:8],2'b0})+$signed(in[583-:8])+$signed({in[591-:8],2'b0})+$signed(in[1039-:8]);
assign sharing20 = $signed({in[615-:8],2'b0})+$signed(in[615-:8])+$signed({in[623-:8],2'b0})+$signed(in[1071-:8]);
assign sharing21 = $signed({in[631-:8],2'b0})+$signed(in[631-:8])+$signed({in[639-:8],2'b0})+$signed(in[1087-:8]);
assign sharing22 = $signed({in[647-:8],2'b0})+$signed(in[647-:8])+$signed({in[655-:8],2'b0})+$signed(in[1103-:8]);
assign sharing23 = $signed({in[903-:8],2'b0})+$signed(in[903-:8])+$signed({in[911-:8],2'b0})+$signed(in[1359-:8]);
assign sharing24 = $signed({in[919-:8],2'b0})+$signed(in[919-:8])+$signed({in[927-:8],2'b0})+$signed(in[1375-:8]);
assign sharing25 = $signed({in[935-:8],2'b0})+$signed(in[935-:8])+$signed({in[943-:8],2'b0})+$signed(in[1391-:8]);
assign sharing26 = $signed({in[951-:8],2'b0})+$signed(in[951-:8])+$signed({in[959-:8],2'b0})+$signed(in[1407-:8]);
assign sharing27 = $signed({in[983-:8],2'b0})+$signed(in[983-:8])+$signed({in[991-:8],2'b0})+$signed(in[1439-:8]);
assign sharing28 = $signed({in[999-:8],2'b0})+$signed(in[999-:8])+$signed({in[1007-:8],2'b0})+$signed(in[1455-:8]);
assign sharing29 = $signed({in[1015-:8],2'b0})+$signed(in[1015-:8])+$signed({in[1023-:8],2'b0})+$signed(in[1471-:8]);
assign sharing30 = $signed({in[1031-:8],2'b0})+$signed(in[1031-:8])+$signed({in[1039-:8],2'b0})+$signed(in[1487-:8]);
assign sharing31 = $signed({in[1047-:8],2'b0})+$signed(in[1047-:8])+$signed({in[1055-:8],2'b0})+$signed(in[1503-:8]);
assign sharing32 = $signed({in[1063-:8],2'b0})+$signed(in[1063-:8])+$signed({in[1071-:8],2'b0})+$signed(in[1519-:8]);
assign sharing33 = $signed({in[1079-:8],2'b0})+$signed(in[1079-:8])+$signed({in[1087-:8],2'b0})+$signed(in[1535-:8]);
assign sharing34 = $signed({in[1351-:8],2'b0})+$signed(in[1351-:8])+$signed({in[1359-:8],2'b0})+$signed(in[1807-:8]);
assign sharing35 = $signed({in[1367-:8],2'b0})+$signed(in[1367-:8])+$signed({in[1375-:8],2'b0})+$signed(in[1823-:8]);
assign sharing36 = $signed({in[1383-:8],2'b0})+$signed(in[1383-:8])+$signed({in[1391-:8],2'b0})+$signed(in[1839-:8]);
assign sharing37 = $signed({in[1399-:8],2'b0})+$signed(in[1399-:8])+$signed({in[1407-:8],2'b0})+$signed(in[1855-:8]);
assign sharing38 = $signed({in[1415-:8],2'b0})+$signed(in[1415-:8])+$signed({in[1423-:8],2'b0})+$signed(in[1871-:8]);
assign sharing39 = $signed({in[1431-:8],2'b0})+$signed(in[1431-:8])+$signed({in[1439-:8],2'b0})+$signed(in[1887-:8]);
assign sharing40 = $signed({in[1447-:8],2'b0})+$signed(in[1447-:8])+$signed({in[1455-:8],2'b0})+$signed(in[1903-:8]);
assign sharing41 = $signed({in[1479-:8],2'b0})+$signed(in[1479-:8])+$signed({in[1487-:8],2'b0})+$signed(in[1935-:8]);
assign sharing42 = $signed({in[1495-:8],2'b0})+$signed(in[1495-:8])+$signed({in[1503-:8],2'b0})+$signed(in[1951-:8]);
assign sharing43 = $signed({in[1511-:8],2'b0})+$signed(in[1511-:8])+$signed({in[1519-:8],2'b0})+$signed(in[1967-:8]);
assign sharing44 = $signed({in[1527-:8],2'b0})+$signed(in[1527-:8])+$signed({in[1535-:8],2'b0})+$signed(in[1983-:8]);
assign sharing45 = $signed({in[1543-:8],2'b0})+$signed(in[1543-:8])+$signed({in[1551-:8],2'b0})+$signed(in[1999-:8]);
assign sharing46 = $signed({in[1799-:8],2'b0})+$signed(in[1799-:8])+$signed({in[1807-:8],2'b0})+$signed(in[2255-:8]);
assign sharing47 = $signed({in[1815-:8],2'b0})+$signed(in[1815-:8])+$signed({in[1823-:8],2'b0})+$signed(in[2271-:8]);
assign sharing48 = $signed({in[1847-:8],2'b0})+$signed(in[1847-:8])+$signed({in[1855-:8],2'b0})+$signed(in[2303-:8]);
assign sharing49 = $signed({in[1863-:8],2'b0})+$signed(in[1863-:8])+$signed({in[1871-:8],2'b0})+$signed(in[2319-:8]);
assign sharing50 = $signed({in[1879-:8],2'b0})+$signed(in[1879-:8])+$signed({in[1887-:8],2'b0})+$signed(in[2335-:8]);
assign sharing51 = $signed({in[1895-:8],2'b0})+$signed(in[1895-:8])+$signed({in[1903-:8],2'b0})+$signed(in[2351-:8]);
assign sharing52 = $signed({in[1911-:8],2'b0})+$signed(in[1911-:8])+$signed({in[1919-:8],2'b0})+$signed(in[2367-:8]);
assign sharing53 = $signed({in[1927-:8],2'b0})+$signed(in[1927-:8])+$signed({in[1935-:8],2'b0})+$signed(in[2383-:8]);
assign sharing54 = $signed({in[1943-:8],2'b0})+$signed(in[1943-:8])+$signed({in[1951-:8],2'b0})+$signed(in[2399-:8]);
assign sharing55 = $signed({in[1975-:8],2'b0})+$signed(in[1975-:8])+$signed({in[1983-:8],2'b0})+$signed(in[2431-:8]);
assign sharing56 = $signed({in[1991-:8],2'b0})+$signed(in[1991-:8])+$signed({in[1999-:8],2'b0})+$signed(in[2447-:8]);
assign sharing57 = $signed({in[2247-:8],2'b0})+$signed(in[2247-:8])+$signed({in[2255-:8],2'b0})+$signed(in[2703-:8]);
assign sharing58 = $signed({in[2263-:8],2'b0})+$signed(in[2263-:8])+$signed({in[2271-:8],2'b0})+$signed(in[2719-:8]);
assign sharing59 = $signed({in[2279-:8],2'b0})+$signed(in[2279-:8])+$signed({in[2287-:8],2'b0})+$signed(in[2735-:8]);
assign sharing60 = $signed({in[2295-:8],2'b0})+$signed(in[2295-:8])+$signed({in[2303-:8],2'b0})+$signed(in[2751-:8]);
assign sharing61 = $signed({in[2311-:8],2'b0})+$signed(in[2311-:8])+$signed({in[2319-:8],2'b0})+$signed(in[2767-:8]);
assign sharing62 = $signed({in[2343-:8],2'b0})+$signed(in[2343-:8])+$signed({in[2351-:8],2'b0})+$signed(in[2799-:8]);
assign sharing63 = $signed({in[2359-:8],2'b0})+$signed(in[2359-:8])+$signed({in[2367-:8],2'b0})+$signed(in[2815-:8]);
assign sharing64 = $signed({in[2375-:8],2'b0})+$signed(in[2375-:8])+$signed({in[2383-:8],2'b0})+$signed(in[2831-:8]);
assign sharing65 = $signed({in[2391-:8],2'b0})+$signed(in[2391-:8])+$signed({in[2399-:8],2'b0})+$signed(in[2847-:8]);
assign sharing66 = $signed({in[2407-:8],2'b0})+$signed(in[2407-:8])+$signed({in[2415-:8],2'b0})+$signed(in[2863-:8]);
assign sharing67 = $signed({in[2423-:8],2'b0})+$signed(in[2423-:8])+$signed({in[2431-:8],2'b0})+$signed(in[2879-:8]);
assign sharing68 = $signed({in[2439-:8],2'b0})+$signed(in[2439-:8])+$signed({in[2447-:8],2'b0})+$signed(in[2895-:8]);
assign sharing69 = $signed({in[2711-:8],2'b0})+$signed(in[2711-:8])+$signed({in[2719-:8],2'b0})+$signed(in[3167-:8]);
assign sharing70 = $signed({in[2727-:8],2'b0})+$signed(in[2727-:8])+$signed({in[2735-:8],2'b0})+$signed(in[3183-:8]);
assign sharing71 = $signed({in[2743-:8],2'b0})+$signed(in[2743-:8])+$signed({in[2751-:8],2'b0})+$signed(in[3199-:8]);
assign sharing72 = $signed({in[2759-:8],2'b0})+$signed(in[2759-:8])+$signed({in[2767-:8],2'b0})+$signed(in[3215-:8]);
assign sharing73 = $signed({in[2775-:8],2'b0})+$signed(in[2775-:8])+$signed({in[2783-:8],2'b0})+$signed(in[3231-:8]);
assign sharing74 = $signed({in[2791-:8],2'b0})+$signed(in[2791-:8])+$signed({in[2799-:8],2'b0})+$signed(in[3247-:8]);
assign sharing75 = $signed({in[2807-:8],2'b0})+$signed(in[2807-:8])+$signed({in[2815-:8],2'b0})+$signed(in[3263-:8]);
assign sharing76 = $signed({in[2839-:8],2'b0})+$signed(in[2839-:8])+$signed({in[2847-:8],2'b0})+$signed(in[3295-:8]);
assign sharing77 = $signed({in[2855-:8],2'b0})+$signed(in[2855-:8])+$signed({in[2863-:8],2'b0})+$signed(in[3311-:8]);
assign sharing78 = $signed({in[2871-:8],2'b0})+$signed(in[2871-:8])+$signed({in[2879-:8],2'b0})+$signed(in[3327-:8]);
assign sharing79 = $signed({in[2887-:8],2'b0})+$signed(in[2887-:8])+$signed({in[2895-:8],2'b0})+$signed(in[3343-:8]);
assign sharing80 = $signed({in[3143-:8],2'b0})+$signed(in[3143-:8])+$signed({in[3151-:8],2'b0})+$signed(in[3599-:8]);
assign sharing81 = $signed({in[3159-:8],2'b0})+$signed(in[3159-:8])+$signed({in[3167-:8],2'b0})+$signed(in[3615-:8]);
assign sharing82 = $signed({in[3175-:8],2'b0})+$signed(in[3175-:8])+$signed({in[3183-:8],2'b0})+$signed(in[3631-:8]);
assign sharing83 = $signed({in[3207-:8],2'b0})+$signed(in[3207-:8])+$signed({in[3215-:8],2'b0})+$signed(in[3663-:8]);
assign sharing84 = $signed({in[3223-:8],2'b0})+$signed(in[3223-:8])+$signed({in[3231-:8],2'b0})+$signed(in[3679-:8]);
assign sharing85 = $signed({in[3239-:8],2'b0})+$signed(in[3239-:8])+$signed({in[3247-:8],2'b0})+$signed(in[3695-:8]);
assign sharing86 = $signed({in[3255-:8],2'b0})+$signed(in[3255-:8])+$signed({in[3263-:8],2'b0})+$signed(in[3711-:8]);
assign sharing87 = $signed({in[3271-:8],2'b0})+$signed(in[3271-:8])+$signed({in[3279-:8],2'b0})+$signed(in[3727-:8]);
assign sharing88 = $signed({in[3287-:8],2'b0})+$signed(in[3287-:8])+$signed({in[3295-:8],2'b0})+$signed(in[3743-:8]);
assign sharing89 = $signed({in[3303-:8],2'b0})+$signed(in[3303-:8])+$signed({in[3311-:8],2'b0})+$signed(in[3759-:8]);
assign sharing90 = $signed({in[3335-:8],2'b0})+$signed(in[3335-:8])+$signed({in[3343-:8],2'b0})+$signed(in[3791-:8]);
assign sharing91 = $signed({in[3591-:8],2'b0})+$signed(in[3591-:8])+$signed({in[3599-:8],2'b0})+$signed(in[4047-:8]);
assign sharing92 = $signed({in[3607-:8],2'b0})+$signed(in[3607-:8])+$signed({in[3615-:8],2'b0})+$signed(in[4063-:8]);
assign sharing93 = $signed({in[3623-:8],2'b0})+$signed(in[3623-:8])+$signed({in[3631-:8],2'b0})+$signed(in[4079-:8]);
assign sharing94 = $signed({in[3639-:8],2'b0})+$signed(in[3639-:8])+$signed({in[3647-:8],2'b0})+$signed(in[4095-:8]);
assign sharing95 = $signed({in[3655-:8],2'b0})+$signed(in[3655-:8])+$signed({in[3663-:8],2'b0})+$signed(in[4111-:8]);
assign sharing96 = $signed({in[3671-:8],2'b0})+$signed(in[3671-:8])+$signed({in[3679-:8],2'b0})+$signed(in[4127-:8]);
assign sharing97 = $signed({in[3703-:8],2'b0})+$signed(in[3703-:8])+$signed({in[3711-:8],2'b0})+$signed(in[4159-:8]);
assign sharing98 = $signed({in[3719-:8],2'b0})+$signed(in[3719-:8])+$signed({in[3727-:8],2'b0})+$signed(in[4175-:8]);
assign sharing99 = $signed({in[3735-:8],2'b0})+$signed(in[3735-:8])+$signed({in[3743-:8],2'b0})+$signed(in[4191-:8]);
assign sharing100 = $signed({in[3751-:8],2'b0})+$signed(in[3751-:8])+$signed({in[3759-:8],2'b0})+$signed(in[4207-:8]);
assign sharing101 = $signed({in[3767-:8],2'b0})+$signed(in[3767-:8])+$signed({in[3775-:8],2'b0})+$signed(in[4223-:8]);
assign sharing102 = $signed({in[3783-:8],2'b0})+$signed(in[3783-:8])+$signed({in[3791-:8],2'b0})+$signed(in[4239-:8]);
assign sharing103 = $signed({in[4039-:8],2'b0})+$signed(in[4039-:8])+$signed({in[4047-:8],2'b0})+$signed(in[4495-:8]);
assign sharing104 = $signed({in[4071-:8],2'b0})+$signed(in[4071-:8])+$signed({in[4079-:8],2'b0})+$signed(in[4527-:8]);
assign sharing105 = $signed({in[4087-:8],2'b0})+$signed(in[4087-:8])+$signed({in[4095-:8],2'b0})+$signed(in[4543-:8]);
assign sharing106 = $signed({in[4103-:8],2'b0})+$signed(in[4103-:8])+$signed({in[4111-:8],2'b0})+$signed(in[4559-:8]);
assign sharing107 = $signed({in[4119-:8],2'b0})+$signed(in[4119-:8])+$signed({in[4127-:8],2'b0})+$signed(in[4575-:8]);
assign sharing108 = $signed({in[4135-:8],2'b0})+$signed(in[4135-:8])+$signed({in[4143-:8],2'b0})+$signed(in[4591-:8]);
assign sharing109 = $signed({in[4151-:8],2'b0})+$signed(in[4151-:8])+$signed({in[4159-:8],2'b0})+$signed(in[4607-:8]);
assign sharing110 = $signed({in[4167-:8],2'b0})+$signed(in[4167-:8])+$signed({in[4175-:8],2'b0})+$signed(in[4623-:8]);
assign sharing111 = $signed({in[4199-:8],2'b0})+$signed(in[4199-:8])+$signed({in[4207-:8],2'b0})+$signed(in[4655-:8]);
assign sharing112 = $signed({in[4215-:8],2'b0})+$signed(in[4215-:8])+$signed({in[4223-:8],2'b0})+$signed(in[4671-:8]);
assign sharing113 = $signed({in[4231-:8],2'b0})+$signed(in[4231-:8])+$signed({in[4239-:8],2'b0})+$signed(in[4687-:8]);
assign sharing114 = $signed({in[4487-:8],2'b0})+$signed(in[4487-:8])+$signed({in[4495-:8],2'b0})+$signed(in[4943-:8]);
assign sharing115 = $signed({in[4503-:8],2'b0})+$signed(in[4503-:8])+$signed({in[4511-:8],2'b0})+$signed(in[4959-:8]);
assign sharing116 = $signed({in[4519-:8],2'b0})+$signed(in[4519-:8])+$signed({in[4527-:8],2'b0})+$signed(in[4975-:8]);
assign sharing117 = $signed({in[4535-:8],2'b0})+$signed(in[4535-:8])+$signed({in[4543-:8],2'b0})+$signed(in[4991-:8]);
assign sharing118 = $signed({in[4567-:8],2'b0})+$signed(in[4567-:8])+$signed({in[4575-:8],2'b0})+$signed(in[5023-:8]);
assign sharing119 = $signed({in[4583-:8],2'b0})+$signed(in[4583-:8])+$signed({in[4591-:8],2'b0})+$signed(in[5039-:8]);
assign sharing120 = $signed({in[4599-:8],2'b0})+$signed(in[4599-:8])+$signed({in[4607-:8],2'b0})+$signed(in[5055-:8]);
assign sharing121 = $signed({in[4615-:8],2'b0})+$signed(in[4615-:8])+$signed({in[4623-:8],2'b0})+$signed(in[5071-:8]);
assign sharing122 = $signed({in[4631-:8],2'b0})+$signed(in[4631-:8])+$signed({in[4639-:8],2'b0})+$signed(in[5087-:8]);
assign sharing123 = $signed({in[4647-:8],2'b0})+$signed(in[4647-:8])+$signed({in[4655-:8],2'b0})+$signed(in[5103-:8]);
assign sharing124 = $signed({in[4663-:8],2'b0})+$signed(in[4663-:8])+$signed({in[4671-:8],2'b0})+$signed(in[5119-:8]);
assign sharing125 = $signed({in[4935-:8],2'b0})+$signed(in[4935-:8])+$signed({in[4943-:8],2'b0})+$signed(in[5391-:8]);
assign sharing126 = $signed({in[4951-:8],2'b0})+$signed(in[4951-:8])+$signed({in[4959-:8],2'b0})+$signed(in[5407-:8]);
assign sharing127 = $signed({in[4967-:8],2'b0})+$signed(in[4967-:8])+$signed({in[4975-:8],2'b0})+$signed(in[5423-:8]);
assign sharing128 = $signed({in[4983-:8],2'b0})+$signed(in[4983-:8])+$signed({in[4991-:8],2'b0})+$signed(in[5439-:8]);
assign sharing129 = $signed({in[4999-:8],2'b0})+$signed(in[4999-:8])+$signed({in[5007-:8],2'b0})+$signed(in[5455-:8]);
assign sharing130 = $signed({in[5015-:8],2'b0})+$signed(in[5015-:8])+$signed({in[5023-:8],2'b0})+$signed(in[5471-:8]);
assign sharing131 = $signed({in[5031-:8],2'b0})+$signed(in[5031-:8])+$signed({in[5039-:8],2'b0})+$signed(in[5487-:8]);
assign sharing132 = $signed({in[5063-:8],2'b0})+$signed(in[5063-:8])+$signed({in[5071-:8],2'b0})+$signed(in[5519-:8]);
assign sharing133 = $signed({in[5079-:8],2'b0})+$signed(in[5079-:8])+$signed({in[5087-:8],2'b0})+$signed(in[5535-:8]);
assign sharing134 = $signed({in[5095-:8],2'b0})+$signed(in[5095-:8])+$signed({in[5103-:8],2'b0})+$signed(in[5551-:8]);
assign sharing135 = $signed({in[5111-:8],2'b0})+$signed(in[5111-:8])+$signed({in[5119-:8],2'b0})+$signed(in[5567-:8]);
assign sharing136 = $signed({in[5127-:8],2'b0})+$signed(in[5127-:8])+$signed({in[5135-:8],2'b0})+$signed(in[5583-:8]);
assign sharing137 = $signed({in[5383-:8],2'b0})+$signed(in[5383-:8])+$signed({in[5391-:8],2'b0})+$signed(in[5839-:8]);
assign sharing138 = $signed({in[5399-:8],2'b0})+$signed(in[5399-:8])+$signed({in[5407-:8],2'b0})+$signed(in[5855-:8]);
assign sharing139 = $signed({in[5431-:8],2'b0})+$signed(in[5431-:8])+$signed({in[5439-:8],2'b0})+$signed(in[5887-:8]);
assign sharing140 = $signed({in[5447-:8],2'b0})+$signed(in[5447-:8])+$signed({in[5455-:8],2'b0})+$signed(in[5903-:8]);
assign sharing141 = $signed({in[5463-:8],2'b0})+$signed(in[5463-:8])+$signed({in[5471-:8],2'b0})+$signed(in[5919-:8]);
assign sharing142 = $signed({in[5479-:8],2'b0})+$signed(in[5479-:8])+$signed({in[5487-:8],2'b0})+$signed(in[5935-:8]);
assign sharing143 = $signed({in[5495-:8],2'b0})+$signed(in[5495-:8])+$signed({in[5503-:8],2'b0})+$signed(in[5951-:8]);
assign sharing144 = $signed({in[5511-:8],2'b0})+$signed(in[5511-:8])+$signed({in[5519-:8],2'b0})+$signed(in[5967-:8]);
assign sharing145 = $signed({in[5527-:8],2'b0})+$signed(in[5527-:8])+$signed({in[5535-:8],2'b0})+$signed(in[5983-:8]);
assign sharing146 = $signed({in[5559-:8],2'b0})+$signed(in[5559-:8])+$signed({in[5567-:8],2'b0})+$signed(in[6015-:8]);
assign sharing147 = $signed({in[5575-:8],2'b0})+$signed(in[5575-:8])+$signed({in[5583-:8],2'b0})+$signed(in[6031-:8]);
assign sharing148 = $signed({in[103-:8],2'b0})+$signed(in[103-:8])+$signed({in[111-:8],2'b0})+$signed(in[559-:8]);
assign sharing149 = $signed({in[471-:8],2'b0})+$signed(in[471-:8])+$signed({in[479-:8],2'b0})+$signed(in[927-:8]);
assign sharing150 = $signed({in[599-:8],2'b0})+$signed(in[599-:8])+$signed({in[607-:8],2'b0})+$signed(in[1055-:8]);
assign sharing151 = $signed({in[967-:8],2'b0})+$signed(in[967-:8])+$signed({in[975-:8],2'b0})+$signed(in[1423-:8]);
assign sharing152 = $signed({in[1095-:8],2'b0})+$signed(in[1095-:8])+$signed({in[1103-:8],2'b0})+$signed(in[1551-:8]);
assign sharing153 = $signed({in[1463-:8],2'b0})+$signed(in[1463-:8])+$signed({in[1471-:8],2'b0})+$signed(in[1919-:8]);
assign sharing154 = $signed({in[1831-:8],2'b0})+$signed(in[1831-:8])+$signed({in[1839-:8],2'b0})+$signed(in[2287-:8]);
assign sharing155 = $signed({in[1959-:8],2'b0})+$signed(in[1959-:8])+$signed({in[1967-:8],2'b0})+$signed(in[2415-:8]);
assign sharing156 = $signed({in[2327-:8],2'b0})+$signed(in[2327-:8])+$signed({in[2335-:8],2'b0})+$signed(in[2783-:8]);
assign sharing157 = $signed({in[2695-:8],2'b0})+$signed(in[2695-:8])+$signed({in[2703-:8],2'b0})+$signed(in[3151-:8]);
assign sharing158 = $signed({in[2823-:8],2'b0})+$signed(in[2823-:8])+$signed({in[2831-:8],2'b0})+$signed(in[3279-:8]);
assign sharing159 = $signed({in[3191-:8],2'b0})+$signed(in[3191-:8])+$signed({in[3199-:8],2'b0})+$signed(in[3647-:8]);
assign sharing160 = $signed({in[3319-:8],2'b0})+$signed(in[3319-:8])+$signed({in[3327-:8],2'b0})+$signed(in[3775-:8]);
assign sharing161 = $signed({in[3687-:8],2'b0})+$signed(in[3687-:8])+$signed({in[3695-:8],2'b0})+$signed(in[4143-:8]);
assign sharing162 = $signed({in[4055-:8],2'b0})+$signed(in[4055-:8])+$signed({in[4063-:8],2'b0})+$signed(in[4511-:8]);
assign sharing163 = $signed({in[4183-:8],2'b0})+$signed(in[4183-:8])+$signed({in[4191-:8],2'b0})+$signed(in[4639-:8]);
assign sharing164 = $signed({in[4551-:8],2'b0})+$signed(in[4551-:8])+$signed({in[4559-:8],2'b0})+$signed(in[5007-:8]);
assign sharing165 = $signed({in[4679-:8],2'b0})+$signed(in[4679-:8])+$signed({in[4687-:8],2'b0})+$signed(in[5135-:8]);
assign sharing166 = $signed({in[5047-:8],2'b0})+$signed(in[5047-:8])+$signed({in[5055-:8],2'b0})+$signed(in[5503-:8]);
assign sharing167 = $signed({in[5415-:8],2'b0})+$signed(in[5415-:8])+$signed({in[5423-:8],2'b0})+$signed(in[5871-:8]);
assign sharing168 = $signed({in[5543-:8],2'b0})+$signed(in[5543-:8])+$signed({in[5551-:8],2'b0})+$signed(in[5999-:8]);
assign weighted_sum[0] = $signed(in[7-:8])+$signed(-in[455-:8])+$signed(in[15-:8])+$signed({in[231-:8],2'b0})+$signed(in[231-:8])+$signed({in[239-:8],1'b0})+$signed(in[239-:8])+$signed({in[247-:8],2'b0})+$signed(7);
assign weighted_sum[1] = $signed({in[263-:8],2'b0})+$signed(in[23-:8])+$signed(-in[471-:8])+$signed(in[31-:8])+$signed({in[247-:8],2'b0})+$signed(in[247-:8])+$signed({in[255-:8],1'b0})+$signed(in[255-:8])+$signed(7);
assign weighted_sum[2] = $signed({in[263-:8],2'b0})+$signed(in[263-:8])+$signed({in[271-:8],1'b0})+$signed(in[271-:8])+$signed({in[279-:8],2'b0})+$signed(in[39-:8])+$signed(-in[487-:8])+$signed(in[47-:8])+$signed(7);
assign weighted_sum[3] = $signed(in[55-:8])+$signed({in[279-:8],2'b0})+$signed(in[279-:8])+$signed({in[287-:8],1'b0})+$signed(in[287-:8])+$signed({in[295-:8],2'b0})+$signed(-in[503-:8])+$signed(in[63-:8])+$signed(7);
assign weighted_sum[4] = $signed(-in[519-:8])+$signed(in[71-:8])+$signed(in[79-:8])+$signed({in[295-:8],2'b0})+$signed(in[295-:8])+$signed({in[303-:8],1'b0})+$signed(in[303-:8])+$signed({in[311-:8],2'b0})+$signed(7);
assign weighted_sum[5] = $signed({in[327-:8],2'b0})+$signed(-in[535-:8])+$signed(in[87-:8])+$signed(in[95-:8])+$signed({in[311-:8],2'b0})+$signed(in[311-:8])+$signed({in[319-:8],1'b0})+$signed(in[319-:8])+$signed(7);
assign weighted_sum[6] = $signed({in[327-:8],2'b0})+$signed(in[327-:8])+$signed({in[335-:8],1'b0})+$signed(in[335-:8])+$signed({in[343-:8],2'b0})+$signed(in[103-:8])+$signed(-in[551-:8])+$signed(in[111-:8])+$signed(7);
assign weighted_sum[7] = $signed({in[343-:8],2'b0})+$signed(in[119-:8])+$signed(in[343-:8])+$signed({in[351-:8],1'b0})+$signed(in[351-:8])+$signed({in[359-:8],2'b0})+$signed(-in[567-:8])+$signed(in[127-:8])+$signed(7);
assign weighted_sum[8] = $signed(-in[583-:8])+$signed(in[135-:8])+$signed(in[143-:8])+$signed({in[359-:8],2'b0})+$signed(in[359-:8])+$signed({in[367-:8],1'b0})+$signed(in[367-:8])+$signed({in[375-:8],2'b0})+$signed(7);
assign weighted_sum[9] = $signed({in[391-:8],2'b0})+$signed(in[151-:8])+$signed(-in[599-:8])+$signed(in[159-:8])+$signed({in[375-:8],2'b0})+$signed(in[375-:8])+$signed({in[383-:8],1'b0})+$signed(in[383-:8])+$signed(7);
assign weighted_sum[10] = $signed({in[391-:8],2'b0})+$signed(in[391-:8])+$signed({in[399-:8],1'b0})+$signed(in[399-:8])+$signed({in[407-:8],2'b0})+$signed(in[167-:8])+$signed(-in[615-:8])+$signed(in[175-:8])+$signed(7);
assign weighted_sum[11] = $signed({in[407-:8],2'b0})+$signed(in[183-:8])+$signed(in[407-:8])+$signed({in[415-:8],1'b0})+$signed(in[415-:8])+$signed({in[423-:8],2'b0})+$signed(-in[631-:8])+$signed(in[191-:8])+$signed(7);
assign weighted_sum[12] = $signed(-in[647-:8])+$signed(in[199-:8])+$signed(in[207-:8])+$signed({in[423-:8],2'b0})+$signed(in[423-:8])+$signed({in[431-:8],1'b0})+$signed(in[431-:8])+$signed({in[439-:8],2'b0})+$signed(7);
assign weighted_sum[13] = $signed(in[455-:8])+$signed(-in[903-:8])+$signed(in[463-:8])+$signed({in[679-:8],2'b0})+$signed(in[679-:8])+$signed({in[687-:8],1'b0})+$signed(in[687-:8])+$signed({in[695-:8],2'b0})+$signed(7);
assign weighted_sum[14] = $signed({in[711-:8],2'b0})+$signed(in[471-:8])+$signed(-in[919-:8])+$signed(in[479-:8])+$signed({in[695-:8],2'b0})+$signed(in[695-:8])+$signed({in[703-:8],1'b0})+$signed(in[703-:8])+$signed(7);
assign weighted_sum[15] = $signed({in[711-:8],2'b0})+$signed(in[711-:8])+$signed({in[719-:8],1'b0})+$signed(in[719-:8])+$signed({in[727-:8],2'b0})+$signed(in[487-:8])+$signed(-in[935-:8])+$signed(in[495-:8])+$signed(7);
assign weighted_sum[16] = $signed({in[727-:8],2'b0})+$signed(in[727-:8])+$signed({in[735-:8],1'b0})+$signed(in[735-:8])+$signed(in[503-:8])+$signed({in[743-:8],2'b0})+$signed(-in[951-:8])+$signed(in[511-:8])+$signed(7);
assign weighted_sum[17] = $signed(in[519-:8])+$signed(-in[967-:8])+$signed(in[527-:8])+$signed({in[743-:8],2'b0})+$signed(in[743-:8])+$signed({in[751-:8],1'b0})+$signed(in[751-:8])+$signed({in[759-:8],2'b0})+$signed(7);
assign weighted_sum[18] = $signed({in[775-:8],2'b0})+$signed(in[535-:8])+$signed(-in[983-:8])+$signed(in[543-:8])+$signed({in[759-:8],2'b0})+$signed(in[759-:8])+$signed({in[767-:8],1'b0})+$signed(in[767-:8])+$signed(7);
assign weighted_sum[19] = $signed({in[775-:8],2'b0})+$signed(in[775-:8])+$signed({in[783-:8],1'b0})+$signed(in[783-:8])+$signed({in[791-:8],2'b0})+$signed(in[551-:8])+$signed(-in[999-:8])+$signed(in[559-:8])+$signed(7);
assign weighted_sum[20] = $signed({in[791-:8],2'b0})+$signed(in[791-:8])+$signed({in[799-:8],1'b0})+$signed(in[799-:8])+$signed(in[567-:8])+$signed({in[807-:8],2'b0})+$signed(-in[1015-:8])+$signed(in[575-:8])+$signed(7);
assign weighted_sum[21] = $signed(-in[1031-:8])+$signed(in[583-:8])+$signed(in[591-:8])+$signed({in[807-:8],2'b0})+$signed(in[807-:8])+$signed({in[815-:8],1'b0})+$signed(in[815-:8])+$signed({in[823-:8],2'b0})+$signed(7);
assign weighted_sum[22] = $signed({in[839-:8],2'b0})+$signed(-in[1047-:8])+$signed(in[599-:8])+$signed(in[607-:8])+$signed({in[823-:8],2'b0})+$signed(in[823-:8])+$signed({in[831-:8],1'b0})+$signed(in[831-:8])+$signed(7);
assign weighted_sum[23] = $signed({in[839-:8],2'b0})+$signed(in[839-:8])+$signed({in[847-:8],1'b0})+$signed(in[847-:8])+$signed({in[855-:8],2'b0})+$signed(in[615-:8])+$signed(-in[1063-:8])+$signed(in[623-:8])+$signed(7);
assign weighted_sum[24] = $signed({in[855-:8],2'b0})+$signed(in[855-:8])+$signed({in[863-:8],1'b0})+$signed(in[863-:8])+$signed({in[871-:8],2'b0})+$signed(in[631-:8])+$signed(-in[1079-:8])+$signed(in[639-:8])+$signed(7);
assign weighted_sum[25] = $signed(-in[1095-:8])+$signed(in[647-:8])+$signed(in[655-:8])+$signed({in[871-:8],2'b0})+$signed(in[871-:8])+$signed({in[879-:8],1'b0})+$signed(in[879-:8])+$signed({in[887-:8],2'b0})+$signed(7);
assign weighted_sum[26] = $signed(in[903-:8])+$signed(-in[1351-:8])+$signed(in[911-:8])+$signed({in[1127-:8],2'b0})+$signed(in[1127-:8])+$signed({in[1135-:8],1'b0})+$signed(in[1135-:8])+$signed({in[1143-:8],2'b0})+$signed(7);
assign weighted_sum[27] = $signed({in[1159-:8],2'b0})+$signed(in[919-:8])+$signed(-in[1367-:8])+$signed(in[927-:8])+$signed({in[1143-:8],2'b0})+$signed(in[1143-:8])+$signed({in[1151-:8],1'b0})+$signed(in[1151-:8])+$signed(7);
assign weighted_sum[28] = $signed({in[1159-:8],2'b0})+$signed(in[1159-:8])+$signed({in[1167-:8],1'b0})+$signed(in[1167-:8])+$signed({in[1175-:8],2'b0})+$signed(in[935-:8])+$signed(-in[1383-:8])+$signed(in[943-:8])+$signed(7);
assign weighted_sum[29] = $signed({in[1175-:8],2'b0})+$signed(in[1175-:8])+$signed({in[1183-:8],1'b0})+$signed(in[1183-:8])+$signed({in[1191-:8],2'b0})+$signed(in[951-:8])+$signed(-in[1399-:8])+$signed(in[959-:8])+$signed(7);
assign weighted_sum[30] = $signed(in[967-:8])+$signed(-in[1415-:8])+$signed(in[975-:8])+$signed({in[1191-:8],2'b0})+$signed(in[1191-:8])+$signed({in[1199-:8],1'b0})+$signed(in[1199-:8])+$signed({in[1207-:8],2'b0})+$signed(7);
assign weighted_sum[31] = $signed({in[1223-:8],2'b0})+$signed(in[983-:8])+$signed(-in[1431-:8])+$signed(in[991-:8])+$signed({in[1207-:8],2'b0})+$signed(in[1207-:8])+$signed({in[1215-:8],1'b0})+$signed(in[1215-:8])+$signed(7);
assign weighted_sum[32] = $signed({in[1223-:8],2'b0})+$signed(in[1223-:8])+$signed({in[1231-:8],1'b0})+$signed(in[1231-:8])+$signed({in[1239-:8],2'b0})+$signed(in[999-:8])+$signed(-in[1447-:8])+$signed(in[1007-:8])+$signed(7);
assign weighted_sum[33] = $signed({in[1239-:8],2'b0})+$signed(in[1239-:8])+$signed({in[1247-:8],1'b0})+$signed(in[1247-:8])+$signed({in[1255-:8],2'b0})+$signed(in[1015-:8])+$signed(-in[1463-:8])+$signed(in[1023-:8])+$signed(7);
assign weighted_sum[34] = $signed(in[1031-:8])+$signed(-in[1479-:8])+$signed(in[1039-:8])+$signed({in[1255-:8],2'b0})+$signed(in[1255-:8])+$signed({in[1263-:8],1'b0})+$signed(in[1263-:8])+$signed({in[1271-:8],2'b0})+$signed(7);
assign weighted_sum[35] = $signed({in[1287-:8],2'b0})+$signed(in[1047-:8])+$signed(-in[1495-:8])+$signed(in[1055-:8])+$signed({in[1271-:8],2'b0})+$signed(in[1271-:8])+$signed({in[1279-:8],1'b0})+$signed(in[1279-:8])+$signed(7);
assign weighted_sum[36] = $signed({in[1287-:8],2'b0})+$signed(in[1287-:8])+$signed({in[1295-:8],1'b0})+$signed(in[1295-:8])+$signed({in[1303-:8],2'b0})+$signed(in[1063-:8])+$signed(-in[1511-:8])+$signed(in[1071-:8])+$signed(7);
assign weighted_sum[37] = $signed({in[1303-:8],2'b0})+$signed(in[1303-:8])+$signed(in[1087-:8])+$signed({in[1311-:8],1'b0})+$signed(in[1311-:8])+$signed({in[1319-:8],2'b0})+$signed(in[1079-:8])+$signed(-in[1527-:8])+$signed(7);
assign weighted_sum[38] = $signed(-in[1543-:8])+$signed(in[1095-:8])+$signed(in[1103-:8])+$signed({in[1319-:8],2'b0})+$signed(in[1319-:8])+$signed({in[1327-:8],1'b0})+$signed(in[1327-:8])+$signed({in[1335-:8],2'b0})+$signed(7);
assign weighted_sum[39] = $signed(in[1351-:8])+$signed(-in[1799-:8])+$signed(in[1359-:8])+$signed({in[1575-:8],2'b0})+$signed(in[1575-:8])+$signed({in[1583-:8],1'b0})+$signed(in[1583-:8])+$signed({in[1591-:8],2'b0})+$signed(7);
assign weighted_sum[40] = $signed({in[1607-:8],2'b0})+$signed(in[1367-:8])+$signed(-in[1815-:8])+$signed(in[1375-:8])+$signed({in[1591-:8],2'b0})+$signed(in[1591-:8])+$signed({in[1599-:8],1'b0})+$signed(in[1599-:8])+$signed(7);
assign weighted_sum[41] = $signed({in[1607-:8],2'b0})+$signed(in[1607-:8])+$signed({in[1615-:8],1'b0})+$signed(in[1615-:8])+$signed({in[1623-:8],2'b0})+$signed(in[1383-:8])+$signed(-in[1831-:8])+$signed(in[1391-:8])+$signed(7);
assign weighted_sum[42] = $signed({in[1623-:8],2'b0})+$signed(in[1623-:8])+$signed({in[1631-:8],1'b0})+$signed(in[1631-:8])+$signed({in[1639-:8],2'b0})+$signed(-in[1847-:8])+$signed(in[1399-:8])+$signed(in[1407-:8])+$signed(7);
assign weighted_sum[43] = $signed(in[1415-:8])+$signed(-in[1863-:8])+$signed(in[1423-:8])+$signed({in[1639-:8],2'b0})+$signed(in[1639-:8])+$signed({in[1647-:8],1'b0})+$signed(in[1647-:8])+$signed({in[1655-:8],2'b0})+$signed(7);
assign weighted_sum[44] = $signed({in[1671-:8],2'b0})+$signed(in[1431-:8])+$signed(-in[1879-:8])+$signed(in[1439-:8])+$signed({in[1655-:8],2'b0})+$signed(in[1655-:8])+$signed({in[1663-:8],1'b0})+$signed(in[1663-:8])+$signed(7);
assign weighted_sum[45] = $signed({in[1671-:8],2'b0})+$signed(in[1671-:8])+$signed({in[1679-:8],1'b0})+$signed(in[1679-:8])+$signed({in[1687-:8],2'b0})+$signed(in[1447-:8])+$signed(-in[1895-:8])+$signed(in[1455-:8])+$signed(7);
assign weighted_sum[46] = $signed({in[1687-:8],2'b0})+$signed(in[1687-:8])+$signed({in[1695-:8],1'b0})+$signed(in[1695-:8])+$signed({in[1703-:8],2'b0})+$signed(-in[1911-:8])+$signed(in[1463-:8])+$signed(in[1471-:8])+$signed(7);
assign weighted_sum[47] = $signed(in[1479-:8])+$signed(-in[1927-:8])+$signed(in[1487-:8])+$signed({in[1703-:8],2'b0})+$signed(in[1703-:8])+$signed({in[1711-:8],1'b0})+$signed(in[1711-:8])+$signed({in[1719-:8],2'b0})+$signed(7);
assign weighted_sum[48] = $signed({in[1735-:8],2'b0})+$signed(in[1495-:8])+$signed(-in[1943-:8])+$signed(in[1503-:8])+$signed({in[1719-:8],2'b0})+$signed(in[1719-:8])+$signed({in[1727-:8],1'b0})+$signed(in[1727-:8])+$signed(7);
assign weighted_sum[49] = $signed({in[1735-:8],2'b0})+$signed(in[1735-:8])+$signed({in[1743-:8],1'b0})+$signed(in[1743-:8])+$signed({in[1751-:8],2'b0})+$signed(in[1511-:8])+$signed(-in[1959-:8])+$signed(in[1519-:8])+$signed(7);
assign weighted_sum[50] = $signed({in[1751-:8],2'b0})+$signed(in[1751-:8])+$signed({in[1759-:8],1'b0})+$signed(in[1759-:8])+$signed({in[1767-:8],2'b0})+$signed(in[1535-:8])+$signed(-in[1975-:8])+$signed(in[1527-:8])+$signed(7);
assign weighted_sum[51] = $signed(in[1543-:8])+$signed(-in[1991-:8])+$signed(in[1551-:8])+$signed({in[1767-:8],2'b0})+$signed(in[1767-:8])+$signed({in[1775-:8],1'b0})+$signed(in[1775-:8])+$signed({in[1783-:8],2'b0})+$signed(7);
assign weighted_sum[52] = $signed(-in[2247-:8])+$signed(in[1799-:8])+$signed(in[1807-:8])+$signed({in[2023-:8],2'b0})+$signed(in[2023-:8])+$signed({in[2031-:8],1'b0})+$signed(in[2031-:8])+$signed({in[2039-:8],2'b0})+$signed(7);
assign weighted_sum[53] = $signed({in[2055-:8],2'b0})+$signed(in[1815-:8])+$signed(-in[2263-:8])+$signed(in[1823-:8])+$signed({in[2039-:8],2'b0})+$signed(in[2039-:8])+$signed({in[2047-:8],1'b0})+$signed(in[2047-:8])+$signed(7);
assign weighted_sum[54] = $signed({in[2055-:8],2'b0})+$signed(in[2055-:8])+$signed({in[2063-:8],1'b0})+$signed(in[2063-:8])+$signed({in[2071-:8],2'b0})+$signed(in[1831-:8])+$signed(-in[2279-:8])+$signed(in[1839-:8])+$signed(7);
assign weighted_sum[55] = $signed(in[1847-:8])+$signed({in[2071-:8],2'b0})+$signed(in[2071-:8])+$signed({in[2079-:8],1'b0})+$signed(in[2079-:8])+$signed({in[2087-:8],2'b0})+$signed(-in[2295-:8])+$signed(in[1855-:8])+$signed(7);
assign weighted_sum[56] = $signed(in[1863-:8])+$signed(-in[2311-:8])+$signed(in[1871-:8])+$signed({in[2087-:8],2'b0})+$signed(in[2087-:8])+$signed({in[2095-:8],1'b0})+$signed(in[2095-:8])+$signed({in[2103-:8],2'b0})+$signed(7);
assign weighted_sum[57] = $signed({in[2119-:8],2'b0})+$signed(in[1879-:8])+$signed(-in[2327-:8])+$signed(in[1887-:8])+$signed({in[2103-:8],2'b0})+$signed(in[2103-:8])+$signed({in[2111-:8],1'b0})+$signed(in[2111-:8])+$signed(7);
assign weighted_sum[58] = $signed({in[2119-:8],2'b0})+$signed(in[2119-:8])+$signed({in[2127-:8],1'b0})+$signed(in[2127-:8])+$signed({in[2135-:8],2'b0})+$signed(in[1895-:8])+$signed(-in[2343-:8])+$signed(in[1903-:8])+$signed(7);
assign weighted_sum[59] = $signed(in[1911-:8])+$signed({in[2135-:8],2'b0})+$signed(in[2135-:8])+$signed({in[2143-:8],1'b0})+$signed(in[2143-:8])+$signed({in[2151-:8],2'b0})+$signed(-in[2359-:8])+$signed(in[1919-:8])+$signed(7);
assign weighted_sum[60] = $signed(in[1927-:8])+$signed(-in[2375-:8])+$signed(in[1935-:8])+$signed({in[2151-:8],2'b0})+$signed(in[2151-:8])+$signed({in[2159-:8],1'b0})+$signed(in[2159-:8])+$signed({in[2167-:8],2'b0})+$signed(7);
assign weighted_sum[61] = $signed({in[2183-:8],2'b0})+$signed(in[1943-:8])+$signed(-in[2391-:8])+$signed(in[1951-:8])+$signed({in[2167-:8],2'b0})+$signed(in[2167-:8])+$signed({in[2175-:8],1'b0})+$signed(in[2175-:8])+$signed(7);
assign weighted_sum[62] = $signed({in[2183-:8],2'b0})+$signed(in[2183-:8])+$signed({in[2191-:8],1'b0})+$signed(in[2191-:8])+$signed({in[2199-:8],2'b0})+$signed(in[1959-:8])+$signed(-in[2407-:8])+$signed(in[1967-:8])+$signed(7);
assign weighted_sum[63] = $signed(in[1975-:8])+$signed({in[2199-:8],2'b0})+$signed(in[2199-:8])+$signed({in[2207-:8],1'b0})+$signed(in[2207-:8])+$signed({in[2215-:8],2'b0})+$signed(-in[2423-:8])+$signed(in[1983-:8])+$signed(7);
assign weighted_sum[64] = $signed(in[1991-:8])+$signed(-in[2439-:8])+$signed(in[1999-:8])+$signed({in[2215-:8],2'b0})+$signed(in[2215-:8])+$signed({in[2223-:8],1'b0})+$signed(in[2223-:8])+$signed({in[2231-:8],2'b0})+$signed(7);
assign weighted_sum[65] = $signed(-in[2695-:8])+$signed(in[2247-:8])+$signed(in[2255-:8])+$signed({in[2471-:8],2'b0})+$signed(in[2471-:8])+$signed({in[2479-:8],1'b0})+$signed(in[2479-:8])+$signed({in[2487-:8],2'b0})+$signed(7);
assign weighted_sum[66] = $signed({in[2503-:8],2'b0})+$signed(-in[2711-:8])+$signed(in[2263-:8])+$signed(in[2271-:8])+$signed({in[2487-:8],2'b0})+$signed(in[2487-:8])+$signed({in[2495-:8],1'b0})+$signed(in[2495-:8])+$signed(7);
assign weighted_sum[67] = $signed({in[2503-:8],2'b0})+$signed(in[2503-:8])+$signed({in[2511-:8],1'b0})+$signed(in[2511-:8])+$signed({in[2519-:8],2'b0})+$signed(in[2279-:8])+$signed(-in[2727-:8])+$signed(in[2287-:8])+$signed(7);
assign weighted_sum[68] = $signed({in[2519-:8],2'b0})+$signed(in[2519-:8])+$signed(in[2295-:8])+$signed({in[2527-:8],1'b0})+$signed(in[2527-:8])+$signed({in[2535-:8],2'b0})+$signed(-in[2743-:8])+$signed(in[2303-:8])+$signed(7);
assign weighted_sum[69] = $signed(-in[2759-:8])+$signed(in[2311-:8])+$signed(in[2319-:8])+$signed({in[2535-:8],2'b0})+$signed(in[2535-:8])+$signed({in[2543-:8],1'b0})+$signed(in[2543-:8])+$signed({in[2551-:8],2'b0})+$signed(7);
assign weighted_sum[70] = $signed({in[2567-:8],2'b0})+$signed(in[2327-:8])+$signed(-in[2775-:8])+$signed(in[2335-:8])+$signed({in[2551-:8],2'b0})+$signed(in[2551-:8])+$signed({in[2559-:8],1'b0})+$signed(in[2559-:8])+$signed(7);
assign weighted_sum[71] = $signed({in[2567-:8],2'b0})+$signed(in[2567-:8])+$signed({in[2575-:8],1'b0})+$signed(in[2575-:8])+$signed({in[2583-:8],2'b0})+$signed(in[2343-:8])+$signed(-in[2791-:8])+$signed(in[2351-:8])+$signed(7);
assign weighted_sum[72] = $signed({in[2583-:8],2'b0})+$signed(in[2583-:8])+$signed(in[2359-:8])+$signed({in[2591-:8],1'b0})+$signed(in[2591-:8])+$signed({in[2599-:8],2'b0})+$signed(-in[2807-:8])+$signed(in[2367-:8])+$signed(7);
assign weighted_sum[73] = $signed(in[2375-:8])+$signed(-in[2823-:8])+$signed(in[2383-:8])+$signed({in[2599-:8],2'b0})+$signed(in[2599-:8])+$signed({in[2607-:8],1'b0})+$signed(in[2607-:8])+$signed({in[2615-:8],2'b0})+$signed(7);
assign weighted_sum[74] = $signed({in[2631-:8],2'b0})+$signed(in[2391-:8])+$signed(-in[2839-:8])+$signed(in[2399-:8])+$signed({in[2615-:8],2'b0})+$signed(in[2615-:8])+$signed({in[2623-:8],1'b0})+$signed(in[2623-:8])+$signed(7);
assign weighted_sum[75] = $signed({in[2631-:8],2'b0})+$signed(in[2631-:8])+$signed({in[2639-:8],1'b0})+$signed(in[2639-:8])+$signed({in[2647-:8],2'b0})+$signed(in[2407-:8])+$signed(-in[2855-:8])+$signed(in[2415-:8])+$signed(7);
assign weighted_sum[76] = $signed({in[2647-:8],2'b0})+$signed(in[2647-:8])+$signed(in[2423-:8])+$signed({in[2655-:8],1'b0})+$signed(in[2655-:8])+$signed({in[2663-:8],2'b0})+$signed(-in[2871-:8])+$signed(in[2431-:8])+$signed(7);
assign weighted_sum[77] = $signed(in[2439-:8])+$signed(-in[2887-:8])+$signed(in[2447-:8])+$signed({in[2663-:8],2'b0})+$signed(in[2663-:8])+$signed({in[2671-:8],1'b0})+$signed(in[2671-:8])+$signed({in[2679-:8],2'b0})+$signed(7);
assign weighted_sum[78] = $signed(-in[3143-:8])+$signed(in[2695-:8])+$signed(in[2703-:8])+$signed({in[2919-:8],2'b0})+$signed(in[2919-:8])+$signed({in[2927-:8],1'b0})+$signed(in[2927-:8])+$signed({in[2935-:8],2'b0})+$signed(7);
assign weighted_sum[79] = $signed({in[2951-:8],2'b0})+$signed(in[2711-:8])+$signed(-in[3159-:8])+$signed(in[2719-:8])+$signed({in[2935-:8],2'b0})+$signed(in[2935-:8])+$signed({in[2943-:8],1'b0})+$signed(in[2943-:8])+$signed(7);
assign weighted_sum[80] = $signed({in[2951-:8],2'b0})+$signed(in[2951-:8])+$signed({in[2959-:8],1'b0})+$signed(in[2959-:8])+$signed({in[2967-:8],2'b0})+$signed(in[2727-:8])+$signed(-in[3175-:8])+$signed(in[2735-:8])+$signed(7);
assign weighted_sum[81] = $signed({in[2967-:8],2'b0})+$signed(in[2967-:8])+$signed({in[2975-:8],1'b0})+$signed(in[2975-:8])+$signed({in[2983-:8],2'b0})+$signed(in[2743-:8])+$signed(-in[3191-:8])+$signed(in[2751-:8])+$signed(7);
assign weighted_sum[82] = $signed(-in[3207-:8])+$signed(in[2759-:8])+$signed(in[2767-:8])+$signed({in[2983-:8],2'b0})+$signed(in[2983-:8])+$signed({in[2991-:8],1'b0})+$signed(in[2991-:8])+$signed({in[2999-:8],2'b0})+$signed(7);
assign weighted_sum[83] = $signed({in[3015-:8],2'b0})+$signed(-in[3223-:8])+$signed(in[2775-:8])+$signed(in[2783-:8])+$signed({in[2999-:8],2'b0})+$signed(in[2999-:8])+$signed({in[3007-:8],1'b0})+$signed(in[3007-:8])+$signed(7);
assign weighted_sum[84] = $signed({in[3015-:8],2'b0})+$signed(in[3015-:8])+$signed({in[3023-:8],1'b0})+$signed(in[3023-:8])+$signed({in[3031-:8],2'b0})+$signed(in[2791-:8])+$signed(-in[3239-:8])+$signed(in[2799-:8])+$signed(7);
assign weighted_sum[85] = $signed({in[3031-:8],2'b0})+$signed(in[3031-:8])+$signed({in[3039-:8],1'b0})+$signed(in[3039-:8])+$signed({in[3047-:8],2'b0})+$signed(in[2807-:8])+$signed(-in[3255-:8])+$signed(in[2815-:8])+$signed(7);
assign weighted_sum[86] = $signed(-in[3271-:8])+$signed(in[2823-:8])+$signed(in[2831-:8])+$signed({in[3047-:8],2'b0})+$signed(in[3047-:8])+$signed({in[3055-:8],1'b0})+$signed(in[3055-:8])+$signed({in[3063-:8],2'b0})+$signed(7);
assign weighted_sum[87] = $signed({in[3079-:8],2'b0})+$signed(in[2839-:8])+$signed(-in[3287-:8])+$signed(in[2847-:8])+$signed({in[3063-:8],2'b0})+$signed(in[3063-:8])+$signed({in[3071-:8],1'b0})+$signed(in[3071-:8])+$signed(7);
assign weighted_sum[88] = $signed({in[3079-:8],2'b0})+$signed(in[3079-:8])+$signed({in[3087-:8],1'b0})+$signed(in[3087-:8])+$signed({in[3095-:8],2'b0})+$signed(in[2855-:8])+$signed(-in[3303-:8])+$signed(in[2863-:8])+$signed(7);
assign weighted_sum[89] = $signed({in[3095-:8],2'b0})+$signed(in[3095-:8])+$signed({in[3103-:8],1'b0})+$signed(in[3103-:8])+$signed({in[3111-:8],2'b0})+$signed(in[2871-:8])+$signed(-in[3319-:8])+$signed(in[2879-:8])+$signed(7);
assign weighted_sum[90] = $signed(in[2887-:8])+$signed(-in[3335-:8])+$signed(in[2895-:8])+$signed({in[3111-:8],2'b0})+$signed(in[3111-:8])+$signed({in[3119-:8],1'b0})+$signed(in[3119-:8])+$signed({in[3127-:8],2'b0})+$signed(7);
assign weighted_sum[91] = $signed(-in[3591-:8])+$signed(in[3143-:8])+$signed(in[3151-:8])+$signed({in[3367-:8],2'b0})+$signed(in[3367-:8])+$signed({in[3375-:8],1'b0})+$signed(in[3375-:8])+$signed({in[3383-:8],2'b0})+$signed(7);
assign weighted_sum[92] = $signed({in[3399-:8],2'b0})+$signed(-in[3607-:8])+$signed(in[3159-:8])+$signed(in[3167-:8])+$signed({in[3383-:8],2'b0})+$signed(in[3383-:8])+$signed({in[3391-:8],1'b0})+$signed(in[3391-:8])+$signed(7);
assign weighted_sum[93] = $signed({in[3399-:8],2'b0})+$signed(in[3399-:8])+$signed({in[3407-:8],1'b0})+$signed(in[3407-:8])+$signed({in[3415-:8],2'b0})+$signed(in[3175-:8])+$signed(-in[3623-:8])+$signed(in[3183-:8])+$signed(7);
assign weighted_sum[94] = $signed({in[3415-:8],2'b0})+$signed(in[3415-:8])+$signed({in[3423-:8],1'b0})+$signed(in[3423-:8])+$signed({in[3431-:8],2'b0})+$signed(in[3191-:8])+$signed(-in[3639-:8])+$signed(in[3199-:8])+$signed(7);
assign weighted_sum[95] = $signed(-in[3655-:8])+$signed(in[3207-:8])+$signed(in[3215-:8])+$signed({in[3431-:8],2'b0})+$signed(in[3431-:8])+$signed({in[3439-:8],1'b0})+$signed(in[3439-:8])+$signed({in[3447-:8],2'b0})+$signed(7);
assign weighted_sum[96] = $signed({in[3463-:8],2'b0})+$signed(in[3223-:8])+$signed(-in[3671-:8])+$signed(in[3231-:8])+$signed({in[3447-:8],2'b0})+$signed(in[3447-:8])+$signed({in[3455-:8],1'b0})+$signed(in[3455-:8])+$signed(7);
assign weighted_sum[97] = $signed({in[3463-:8],2'b0})+$signed(in[3463-:8])+$signed({in[3471-:8],1'b0})+$signed(in[3471-:8])+$signed({in[3479-:8],2'b0})+$signed(in[3239-:8])+$signed(-in[3687-:8])+$signed(in[3247-:8])+$signed(7);
assign weighted_sum[98] = $signed({in[3479-:8],2'b0})+$signed(in[3479-:8])+$signed({in[3487-:8],1'b0})+$signed(in[3487-:8])+$signed({in[3495-:8],2'b0})+$signed(in[3255-:8])+$signed(-in[3703-:8])+$signed(in[3263-:8])+$signed(7);
assign weighted_sum[99] = $signed(-in[3719-:8])+$signed(in[3271-:8])+$signed(in[3279-:8])+$signed({in[3495-:8],2'b0})+$signed(in[3495-:8])+$signed({in[3503-:8],1'b0})+$signed(in[3503-:8])+$signed({in[3511-:8],2'b0})+$signed(7);
assign weighted_sum[100] = $signed({in[3527-:8],2'b0})+$signed(-in[3735-:8])+$signed(in[3287-:8])+$signed(in[3295-:8])+$signed({in[3511-:8],2'b0})+$signed(in[3511-:8])+$signed({in[3519-:8],1'b0})+$signed(in[3519-:8])+$signed(7);
assign weighted_sum[101] = $signed({in[3527-:8],2'b0})+$signed(in[3527-:8])+$signed({in[3535-:8],1'b0})+$signed(in[3535-:8])+$signed({in[3543-:8],2'b0})+$signed(in[3303-:8])+$signed(-in[3751-:8])+$signed(in[3311-:8])+$signed(7);
assign weighted_sum[102] = $signed({in[3543-:8],2'b0})+$signed(in[3319-:8])+$signed(in[3543-:8])+$signed({in[3551-:8],1'b0})+$signed(in[3551-:8])+$signed({in[3559-:8],2'b0})+$signed(-in[3767-:8])+$signed(in[3327-:8])+$signed(7);
assign weighted_sum[103] = $signed(-in[3783-:8])+$signed(in[3335-:8])+$signed(in[3343-:8])+$signed({in[3559-:8],2'b0})+$signed(in[3559-:8])+$signed({in[3567-:8],1'b0})+$signed(in[3567-:8])+$signed({in[3575-:8],2'b0})+$signed(7);
assign weighted_sum[104] = $signed(in[3591-:8])+$signed(-in[4039-:8])+$signed(in[3599-:8])+$signed({in[3815-:8],2'b0})+$signed(in[3815-:8])+$signed({in[3823-:8],1'b0})+$signed(in[3823-:8])+$signed({in[3831-:8],2'b0})+$signed(7);
assign weighted_sum[105] = $signed({in[3847-:8],2'b0})+$signed(in[3607-:8])+$signed(-in[4055-:8])+$signed(in[3615-:8])+$signed({in[3831-:8],2'b0})+$signed(in[3831-:8])+$signed({in[3839-:8],1'b0})+$signed(in[3839-:8])+$signed(7);
assign weighted_sum[106] = $signed({in[3847-:8],2'b0})+$signed(in[3847-:8])+$signed({in[3855-:8],1'b0})+$signed(in[3855-:8])+$signed({in[3863-:8],2'b0})+$signed(in[3623-:8])+$signed(-in[4071-:8])+$signed(in[3631-:8])+$signed(7);
assign weighted_sum[107] = $signed(in[3639-:8])+$signed({in[3863-:8],2'b0})+$signed(in[3863-:8])+$signed({in[3871-:8],1'b0})+$signed(in[3871-:8])+$signed({in[3879-:8],2'b0})+$signed(-in[4087-:8])+$signed(in[3647-:8])+$signed(7);
assign weighted_sum[108] = $signed(-in[4103-:8])+$signed(in[3655-:8])+$signed(in[3663-:8])+$signed({in[3879-:8],2'b0})+$signed(in[3879-:8])+$signed({in[3887-:8],1'b0})+$signed(in[3887-:8])+$signed({in[3895-:8],2'b0})+$signed(7);
assign weighted_sum[109] = $signed({in[3911-:8],2'b0})+$signed(-in[4119-:8])+$signed(in[3671-:8])+$signed(in[3679-:8])+$signed({in[3895-:8],2'b0})+$signed(in[3895-:8])+$signed({in[3903-:8],1'b0})+$signed(in[3903-:8])+$signed(7);
assign weighted_sum[110] = $signed({in[3911-:8],2'b0})+$signed(in[3911-:8])+$signed({in[3919-:8],1'b0})+$signed(in[3919-:8])+$signed({in[3927-:8],2'b0})+$signed(in[3687-:8])+$signed(-in[4135-:8])+$signed(in[3695-:8])+$signed(7);
assign weighted_sum[111] = $signed(in[3703-:8])+$signed({in[3927-:8],2'b0})+$signed(in[3927-:8])+$signed({in[3935-:8],1'b0})+$signed(in[3935-:8])+$signed({in[3943-:8],2'b0})+$signed(-in[4151-:8])+$signed(in[3711-:8])+$signed(7);
assign weighted_sum[112] = $signed(-in[4167-:8])+$signed(in[3719-:8])+$signed(in[3727-:8])+$signed({in[3943-:8],2'b0})+$signed(in[3943-:8])+$signed({in[3951-:8],1'b0})+$signed(in[3951-:8])+$signed({in[3959-:8],2'b0})+$signed(7);
assign weighted_sum[113] = $signed({in[3975-:8],2'b0})+$signed(-in[4183-:8])+$signed(in[3735-:8])+$signed(in[3743-:8])+$signed({in[3959-:8],2'b0})+$signed(in[3959-:8])+$signed({in[3967-:8],1'b0})+$signed(in[3967-:8])+$signed(7);
assign weighted_sum[114] = $signed({in[3975-:8],2'b0})+$signed(in[3975-:8])+$signed({in[3983-:8],1'b0})+$signed(in[3983-:8])+$signed({in[3991-:8],2'b0})+$signed(in[3751-:8])+$signed(-in[4199-:8])+$signed(in[3759-:8])+$signed(7);
assign weighted_sum[115] = $signed(in[3767-:8])+$signed({in[3991-:8],2'b0})+$signed(in[3991-:8])+$signed({in[3999-:8],1'b0})+$signed(in[3999-:8])+$signed({in[4007-:8],2'b0})+$signed(-in[4215-:8])+$signed(in[3775-:8])+$signed(7);
assign weighted_sum[116] = $signed(-in[4231-:8])+$signed(in[3783-:8])+$signed(in[3791-:8])+$signed({in[4007-:8],2'b0})+$signed(in[4007-:8])+$signed({in[4015-:8],1'b0})+$signed(in[4015-:8])+$signed({in[4023-:8],2'b0})+$signed(7);
assign weighted_sum[117] = $signed(in[4039-:8])+$signed(-in[4487-:8])+$signed(in[4047-:8])+$signed({in[4263-:8],2'b0})+$signed(in[4263-:8])+$signed({in[4271-:8],1'b0})+$signed(in[4271-:8])+$signed({in[4279-:8],2'b0})+$signed(7);
assign weighted_sum[118] = $signed({in[4295-:8],2'b0})+$signed(in[4055-:8])+$signed(-in[4503-:8])+$signed(in[4063-:8])+$signed({in[4279-:8],2'b0})+$signed(in[4279-:8])+$signed({in[4287-:8],1'b0})+$signed(in[4287-:8])+$signed(7);
assign weighted_sum[119] = $signed({in[4295-:8],2'b0})+$signed(in[4295-:8])+$signed({in[4303-:8],1'b0})+$signed(in[4303-:8])+$signed({in[4311-:8],2'b0})+$signed(in[4071-:8])+$signed(-in[4519-:8])+$signed(in[4079-:8])+$signed(7);
assign weighted_sum[120] = $signed(in[4087-:8])+$signed({in[4311-:8],2'b0})+$signed(in[4311-:8])+$signed({in[4319-:8],1'b0})+$signed(in[4319-:8])+$signed({in[4327-:8],2'b0})+$signed(-in[4535-:8])+$signed(in[4095-:8])+$signed(7);
assign weighted_sum[121] = $signed(in[4103-:8])+$signed(-in[4551-:8])+$signed(in[4111-:8])+$signed({in[4327-:8],2'b0})+$signed(in[4327-:8])+$signed({in[4335-:8],1'b0})+$signed(in[4335-:8])+$signed({in[4343-:8],2'b0})+$signed(7);
assign weighted_sum[122] = $signed({in[4359-:8],2'b0})+$signed(in[4119-:8])+$signed(-in[4567-:8])+$signed(in[4127-:8])+$signed({in[4343-:8],2'b0})+$signed(in[4343-:8])+$signed({in[4351-:8],1'b0})+$signed(in[4351-:8])+$signed(7);
assign weighted_sum[123] = $signed({in[4359-:8],2'b0})+$signed(in[4359-:8])+$signed({in[4367-:8],1'b0})+$signed(in[4367-:8])+$signed({in[4375-:8],2'b0})+$signed(in[4135-:8])+$signed(-in[4583-:8])+$signed(in[4143-:8])+$signed(7);
assign weighted_sum[124] = $signed(in[4151-:8])+$signed({in[4375-:8],2'b0})+$signed(in[4375-:8])+$signed({in[4383-:8],1'b0})+$signed(in[4383-:8])+$signed({in[4391-:8],2'b0})+$signed(-in[4599-:8])+$signed(in[4159-:8])+$signed(7);
assign weighted_sum[125] = $signed(-in[4615-:8])+$signed(in[4167-:8])+$signed(in[4175-:8])+$signed({in[4391-:8],2'b0})+$signed(in[4391-:8])+$signed({in[4399-:8],1'b0})+$signed(in[4399-:8])+$signed({in[4407-:8],2'b0})+$signed(7);
assign weighted_sum[126] = $signed({in[4423-:8],2'b0})+$signed(-in[4631-:8])+$signed(in[4183-:8])+$signed(in[4191-:8])+$signed({in[4407-:8],2'b0})+$signed(in[4407-:8])+$signed({in[4415-:8],1'b0})+$signed(in[4415-:8])+$signed(7);
assign weighted_sum[127] = $signed({in[4423-:8],2'b0})+$signed(in[4423-:8])+$signed({in[4431-:8],1'b0})+$signed(in[4431-:8])+$signed({in[4439-:8],2'b0})+$signed(in[4199-:8])+$signed(-in[4647-:8])+$signed(in[4207-:8])+$signed(7);
assign weighted_sum[128] = $signed({in[4439-:8],2'b0})+$signed(in[4215-:8])+$signed(in[4439-:8])+$signed({in[4447-:8],1'b0})+$signed(in[4447-:8])+$signed({in[4455-:8],2'b0})+$signed(-in[4663-:8])+$signed(in[4223-:8])+$signed(7);
assign weighted_sum[129] = $signed(-in[4679-:8])+$signed(in[4231-:8])+$signed(in[4239-:8])+$signed({in[4455-:8],2'b0})+$signed(in[4455-:8])+$signed({in[4463-:8],1'b0})+$signed(in[4463-:8])+$signed({in[4471-:8],2'b0})+$signed(7);
assign weighted_sum[130] = $signed(in[4487-:8])+$signed(-in[4935-:8])+$signed(in[4495-:8])+$signed({in[4711-:8],2'b0})+$signed(in[4711-:8])+$signed({in[4719-:8],1'b0})+$signed(in[4719-:8])+$signed({in[4727-:8],2'b0})+$signed(7);
assign weighted_sum[131] = $signed({in[4743-:8],2'b0})+$signed(in[4503-:8])+$signed(-in[4951-:8])+$signed(in[4511-:8])+$signed({in[4727-:8],2'b0})+$signed(in[4727-:8])+$signed({in[4735-:8],1'b0})+$signed(in[4735-:8])+$signed(7);
assign weighted_sum[132] = $signed({in[4743-:8],2'b0})+$signed(in[4743-:8])+$signed({in[4751-:8],1'b0})+$signed(in[4751-:8])+$signed({in[4759-:8],2'b0})+$signed(in[4519-:8])+$signed(-in[4967-:8])+$signed(in[4527-:8])+$signed(7);
assign weighted_sum[133] = $signed({in[4759-:8],2'b0})+$signed(in[4759-:8])+$signed({in[4767-:8],1'b0})+$signed(in[4767-:8])+$signed(in[4535-:8])+$signed({in[4775-:8],2'b0})+$signed(-in[4983-:8])+$signed(in[4543-:8])+$signed(7);
assign weighted_sum[134] = $signed(in[4551-:8])+$signed(-in[4999-:8])+$signed(in[4559-:8])+$signed({in[4775-:8],2'b0})+$signed(in[4775-:8])+$signed({in[4783-:8],1'b0})+$signed(in[4783-:8])+$signed({in[4791-:8],2'b0})+$signed(7);
assign weighted_sum[135] = $signed({in[4807-:8],2'b0})+$signed(in[4567-:8])+$signed(-in[5015-:8])+$signed(in[4575-:8])+$signed({in[4791-:8],2'b0})+$signed(in[4791-:8])+$signed({in[4799-:8],1'b0})+$signed(in[4799-:8])+$signed(7);
assign weighted_sum[136] = $signed({in[4807-:8],2'b0})+$signed(in[4807-:8])+$signed({in[4815-:8],1'b0})+$signed(in[4815-:8])+$signed({in[4823-:8],2'b0})+$signed(in[4583-:8])+$signed(-in[5031-:8])+$signed(in[4591-:8])+$signed(7);
assign weighted_sum[137] = $signed({in[4823-:8],2'b0})+$signed(in[4823-:8])+$signed({in[4831-:8],1'b0})+$signed(in[4831-:8])+$signed(in[4599-:8])+$signed({in[4839-:8],2'b0})+$signed(-in[5047-:8])+$signed(in[4607-:8])+$signed(7);
assign weighted_sum[138] = $signed(in[4615-:8])+$signed(-in[5063-:8])+$signed(in[4623-:8])+$signed({in[4839-:8],2'b0})+$signed(in[4839-:8])+$signed({in[4847-:8],1'b0})+$signed(in[4847-:8])+$signed({in[4855-:8],2'b0})+$signed(7);
assign weighted_sum[139] = $signed({in[4871-:8],2'b0})+$signed(in[4631-:8])+$signed(-in[5079-:8])+$signed(in[4639-:8])+$signed({in[4855-:8],2'b0})+$signed(in[4855-:8])+$signed({in[4863-:8],1'b0})+$signed(in[4863-:8])+$signed(7);
assign weighted_sum[140] = $signed({in[4871-:8],2'b0})+$signed(in[4871-:8])+$signed({in[4879-:8],1'b0})+$signed(in[4879-:8])+$signed({in[4887-:8],2'b0})+$signed(in[4647-:8])+$signed(-in[5095-:8])+$signed(in[4655-:8])+$signed(7);
assign weighted_sum[141] = $signed({in[4887-:8],2'b0})+$signed(in[4887-:8])+$signed({in[4895-:8],1'b0})+$signed(in[4895-:8])+$signed(in[4663-:8])+$signed({in[4903-:8],2'b0})+$signed(-in[5111-:8])+$signed(in[4671-:8])+$signed(7);
assign weighted_sum[142] = $signed(-in[5127-:8])+$signed(in[4679-:8])+$signed(in[4687-:8])+$signed({in[4903-:8],2'b0})+$signed(in[4903-:8])+$signed({in[4911-:8],1'b0})+$signed(in[4911-:8])+$signed({in[4919-:8],2'b0})+$signed(7);
assign weighted_sum[143] = $signed(in[4935-:8])+$signed(-in[5383-:8])+$signed(in[4943-:8])+$signed({in[5159-:8],2'b0})+$signed(in[5159-:8])+$signed({in[5167-:8],1'b0})+$signed(in[5167-:8])+$signed({in[5175-:8],2'b0})+$signed(7);
assign weighted_sum[144] = $signed({in[5191-:8],2'b0})+$signed(in[4951-:8])+$signed(-in[5399-:8])+$signed(in[4959-:8])+$signed({in[5175-:8],2'b0})+$signed(in[5175-:8])+$signed({in[5183-:8],1'b0})+$signed(in[5183-:8])+$signed(7);
assign weighted_sum[145] = $signed({in[5191-:8],2'b0})+$signed(in[5191-:8])+$signed({in[5199-:8],1'b0})+$signed(in[5199-:8])+$signed({in[5207-:8],2'b0})+$signed(in[4967-:8])+$signed(-in[5415-:8])+$signed(in[4975-:8])+$signed(7);
assign weighted_sum[146] = $signed({in[5207-:8],2'b0})+$signed(in[5207-:8])+$signed({in[5215-:8],1'b0})+$signed(in[5215-:8])+$signed({in[5223-:8],2'b0})+$signed(in[4983-:8])+$signed(-in[5431-:8])+$signed(in[4991-:8])+$signed(7);
assign weighted_sum[147] = $signed(in[4999-:8])+$signed(-in[5447-:8])+$signed(in[5007-:8])+$signed({in[5223-:8],2'b0})+$signed(in[5223-:8])+$signed({in[5231-:8],1'b0})+$signed(in[5231-:8])+$signed({in[5239-:8],2'b0})+$signed(7);
assign weighted_sum[148] = $signed({in[5255-:8],2'b0})+$signed(in[5015-:8])+$signed(-in[5463-:8])+$signed(in[5023-:8])+$signed({in[5239-:8],2'b0})+$signed(in[5239-:8])+$signed({in[5247-:8],1'b0})+$signed(in[5247-:8])+$signed(7);
assign weighted_sum[149] = $signed({in[5255-:8],2'b0})+$signed(in[5255-:8])+$signed({in[5263-:8],1'b0})+$signed(in[5263-:8])+$signed({in[5271-:8],2'b0})+$signed(in[5031-:8])+$signed(-in[5479-:8])+$signed(in[5039-:8])+$signed(7);
assign weighted_sum[150] = $signed({in[5271-:8],2'b0})+$signed(in[5271-:8])+$signed({in[5279-:8],1'b0})+$signed(in[5279-:8])+$signed({in[5287-:8],2'b0})+$signed(in[5047-:8])+$signed(-in[5495-:8])+$signed(in[5055-:8])+$signed(7);
assign weighted_sum[151] = $signed(in[5063-:8])+$signed(-in[5511-:8])+$signed(in[5071-:8])+$signed({in[5287-:8],2'b0})+$signed(in[5287-:8])+$signed({in[5295-:8],1'b0})+$signed(in[5295-:8])+$signed({in[5303-:8],2'b0})+$signed(7);
assign weighted_sum[152] = $signed({in[5319-:8],2'b0})+$signed(in[5079-:8])+$signed(-in[5527-:8])+$signed(in[5087-:8])+$signed({in[5303-:8],2'b0})+$signed(in[5303-:8])+$signed({in[5311-:8],1'b0})+$signed(in[5311-:8])+$signed(7);
assign weighted_sum[153] = $signed({in[5319-:8],2'b0})+$signed(in[5319-:8])+$signed({in[5327-:8],1'b0})+$signed(in[5327-:8])+$signed({in[5335-:8],2'b0})+$signed(in[5095-:8])+$signed(-in[5543-:8])+$signed(in[5103-:8])+$signed(7);
assign weighted_sum[154] = $signed({in[5335-:8],2'b0})+$signed(in[5335-:8])+$signed({in[5343-:8],1'b0})+$signed(in[5343-:8])+$signed({in[5351-:8],2'b0})+$signed(in[5111-:8])+$signed(-in[5559-:8])+$signed(in[5119-:8])+$signed(7);
assign weighted_sum[155] = $signed(in[5127-:8])+$signed(-in[5575-:8])+$signed(in[5135-:8])+$signed({in[5351-:8],2'b0})+$signed(in[5351-:8])+$signed({in[5359-:8],1'b0})+$signed(in[5359-:8])+$signed({in[5367-:8],2'b0})+$signed(7);
assign weighted_sum[156] = $signed(-in[5831-:8])+$signed(in[5383-:8])+$signed(in[5391-:8])+$signed({in[5607-:8],2'b0})+$signed(in[5607-:8])+$signed({in[5615-:8],1'b0})+$signed(in[5615-:8])+$signed({in[5623-:8],2'b0})+$signed(7);
assign weighted_sum[157] = $signed({in[5639-:8],2'b0})+$signed(-in[5847-:8])+$signed(in[5399-:8])+$signed(in[5407-:8])+$signed({in[5623-:8],2'b0})+$signed(in[5623-:8])+$signed({in[5631-:8],1'b0})+$signed(in[5631-:8])+$signed(7);
assign weighted_sum[158] = $signed({in[5639-:8],2'b0})+$signed(in[5639-:8])+$signed({in[5647-:8],1'b0})+$signed(in[5647-:8])+$signed({in[5655-:8],2'b0})+$signed(in[5415-:8])+$signed(-in[5863-:8])+$signed(in[5423-:8])+$signed(7);
assign weighted_sum[159] = $signed({in[5655-:8],2'b0})+$signed(in[5655-:8])+$signed({in[5663-:8],1'b0})+$signed(in[5663-:8])+$signed({in[5671-:8],2'b0})+$signed(-in[5879-:8])+$signed(in[5431-:8])+$signed(in[5439-:8])+$signed(7);
assign weighted_sum[160] = $signed(in[5447-:8])+$signed(-in[5895-:8])+$signed(in[5455-:8])+$signed({in[5671-:8],2'b0})+$signed(in[5671-:8])+$signed({in[5679-:8],1'b0})+$signed(in[5679-:8])+$signed({in[5687-:8],2'b0})+$signed(7);
assign weighted_sum[161] = $signed({in[5703-:8],2'b0})+$signed(in[5463-:8])+$signed(-in[5911-:8])+$signed(in[5471-:8])+$signed({in[5687-:8],2'b0})+$signed(in[5687-:8])+$signed({in[5695-:8],1'b0})+$signed(in[5695-:8])+$signed(7);
assign weighted_sum[162] = $signed({in[5703-:8],2'b0})+$signed(in[5703-:8])+$signed({in[5711-:8],1'b0})+$signed(in[5711-:8])+$signed({in[5719-:8],2'b0})+$signed(in[5479-:8])+$signed(-in[5927-:8])+$signed(in[5487-:8])+$signed(7);
assign weighted_sum[163] = $signed({in[5719-:8],2'b0})+$signed(in[5719-:8])+$signed({in[5727-:8],1'b0})+$signed(in[5727-:8])+$signed({in[5735-:8],2'b0})+$signed(-in[5943-:8])+$signed(in[5495-:8])+$signed(in[5503-:8])+$signed(7);
assign weighted_sum[164] = $signed(in[5511-:8])+$signed(-in[5959-:8])+$signed(in[5519-:8])+$signed({in[5735-:8],2'b0})+$signed(in[5735-:8])+$signed({in[5743-:8],1'b0})+$signed(in[5743-:8])+$signed({in[5751-:8],2'b0})+$signed(7);
assign weighted_sum[165] = $signed({in[5767-:8],2'b0})+$signed(in[5527-:8])+$signed(-in[5975-:8])+$signed(in[5535-:8])+$signed({in[5751-:8],2'b0})+$signed(in[5751-:8])+$signed({in[5759-:8],1'b0})+$signed(in[5759-:8])+$signed(7);
assign weighted_sum[166] = $signed({in[5767-:8],2'b0})+$signed(in[5767-:8])+$signed({in[5775-:8],1'b0})+$signed(in[5775-:8])+$signed({in[5783-:8],2'b0})+$signed(in[5543-:8])+$signed(-in[5991-:8])+$signed(in[5551-:8])+$signed(7);
assign weighted_sum[167] = $signed({in[5783-:8],2'b0})+$signed(in[5783-:8])+$signed({in[5791-:8],1'b0})+$signed(in[5791-:8])+$signed({in[5799-:8],2'b0})+$signed(-in[6007-:8])+$signed(in[5559-:8])+$signed(in[5567-:8])+$signed(7);
assign weighted_sum[168] = $signed(in[5575-:8])+$signed(-in[6023-:8])+$signed(in[5583-:8])+$signed({in[5799-:8],2'b0})+$signed(in[5799-:8])+$signed({in[5807-:8],1'b0})+$signed(in[5807-:8])+$signed({in[5815-:8],2'b0})+$signed(7);
assign weighted_sum[169] = $signed({in[455-:8],1'b0})+$signed(-{in[463-:8],2'b0})+$signed(-{in[471-:8],2'b0})+$signed(-in[23-:8])+$signed({in[231-:8],1'b0})+$signed(in[231-:8])+$signed(-{in[247-:8],2'b0})+$signed(sharing0)+$signed(1);
assign weighted_sum[170] = $signed(-{in[263-:8],2'b0})+$signed({in[471-:8],1'b0})+$signed(-{in[479-:8],2'b0})+$signed(-{in[487-:8],2'b0})+$signed(-in[39-:8])+$signed({in[247-:8],1'b0})+$signed(in[247-:8])+$signed(sharing1)+$signed(1);
assign weighted_sum[171] = $signed({in[263-:8],1'b0})+$signed(in[263-:8])+$signed(-{in[279-:8],2'b0})+$signed({in[487-:8],1'b0})+$signed(-{in[495-:8],2'b0})+$signed(-{in[503-:8],2'b0})+$signed(-in[55-:8])+$signed(sharing2)+$signed(1);
assign weighted_sum[172] = $signed(-{in[519-:8],2'b0})+$signed(-in[71-:8])+$signed({in[279-:8],1'b0})+$signed(in[279-:8])+$signed(-{in[295-:8],2'b0})+$signed({in[503-:8],1'b0})+$signed(-{in[511-:8],2'b0})+$signed(sharing3)+$signed(1);
assign weighted_sum[173] = $signed({in[519-:8],1'b0})+$signed(-{in[527-:8],2'b0})+$signed(-{in[535-:8],2'b0})+$signed(-in[87-:8])+$signed({in[295-:8],1'b0})+$signed(in[295-:8])+$signed(-{in[311-:8],2'b0})+$signed(sharing4)+$signed(1);
assign weighted_sum[174] = $signed(-{in[327-:8],2'b0})+$signed({in[535-:8],1'b0})+$signed(-{in[543-:8],2'b0})+$signed(-{in[551-:8],2'b0})+$signed(-in[103-:8])+$signed({in[311-:8],1'b0})+$signed(in[311-:8])+$signed(sharing5)+$signed(1);
assign weighted_sum[175] = $signed({in[327-:8],1'b0})+$signed(in[327-:8])+$signed(-{in[343-:8],2'b0})+$signed({in[551-:8],1'b0})+$signed(-{in[559-:8],2'b0})+$signed(-{in[567-:8],2'b0})+$signed(-in[119-:8])+$signed(sharing148)+$signed(1);
assign weighted_sum[176] = $signed(-{in[583-:8],2'b0})+$signed(-in[135-:8])+$signed({in[343-:8],1'b0})+$signed(in[343-:8])+$signed(-{in[359-:8],2'b0})+$signed({in[567-:8],1'b0})+$signed(-{in[575-:8],2'b0})+$signed(sharing6)+$signed(1);
assign weighted_sum[177] = $signed({in[583-:8],1'b0})+$signed(-{in[591-:8],2'b0})+$signed(-{in[599-:8],2'b0})+$signed(-in[151-:8])+$signed({in[359-:8],1'b0})+$signed(in[359-:8])+$signed(-{in[375-:8],2'b0})+$signed(sharing7)+$signed(1);
assign weighted_sum[178] = $signed(-{in[391-:8],2'b0})+$signed({in[599-:8],1'b0})+$signed(-{in[607-:8],2'b0})+$signed(-{in[615-:8],2'b0})+$signed(-in[167-:8])+$signed({in[375-:8],1'b0})+$signed(in[375-:8])+$signed(sharing8)+$signed(1);
assign weighted_sum[179] = $signed({in[391-:8],1'b0})+$signed(in[391-:8])+$signed(-{in[407-:8],2'b0})+$signed({in[615-:8],1'b0})+$signed(-{in[623-:8],2'b0})+$signed(-{in[631-:8],2'b0})+$signed(-in[183-:8])+$signed(sharing9)+$signed(1);
assign weighted_sum[180] = $signed(-{in[647-:8],2'b0})+$signed(-in[199-:8])+$signed({in[407-:8],1'b0})+$signed(in[407-:8])+$signed(-{in[423-:8],2'b0})+$signed({in[631-:8],1'b0})+$signed(-{in[639-:8],2'b0})+$signed(sharing10)+$signed(1);
assign weighted_sum[181] = $signed({in[647-:8],1'b0})+$signed(-{in[655-:8],2'b0})+$signed(-{in[663-:8],2'b0})+$signed(-in[215-:8])+$signed({in[423-:8],1'b0})+$signed(in[423-:8])+$signed(-{in[439-:8],2'b0})+$signed(sharing11)+$signed(1);
assign weighted_sum[182] = $signed({in[903-:8],1'b0})+$signed(-{in[911-:8],2'b0})+$signed(-{in[919-:8],2'b0})+$signed(-in[471-:8])+$signed({in[679-:8],1'b0})+$signed(in[679-:8])+$signed(-{in[695-:8],2'b0})+$signed(sharing12)+$signed(1);
assign weighted_sum[183] = $signed(-{in[711-:8],2'b0})+$signed({in[919-:8],1'b0})+$signed(-{in[927-:8],2'b0})+$signed(-{in[935-:8],2'b0})+$signed(-in[487-:8])+$signed({in[695-:8],1'b0})+$signed(in[695-:8])+$signed(sharing149)+$signed(1);
assign weighted_sum[184] = $signed({in[711-:8],1'b0})+$signed(in[711-:8])+$signed(-{in[727-:8],2'b0})+$signed({in[935-:8],1'b0})+$signed(-{in[943-:8],2'b0})+$signed(-{in[951-:8],2'b0})+$signed(-in[503-:8])+$signed(sharing13)+$signed(1);
assign weighted_sum[185] = $signed(-{in[967-:8],2'b0})+$signed(-in[519-:8])+$signed({in[727-:8],1'b0})+$signed(in[727-:8])+$signed(-{in[743-:8],2'b0})+$signed({in[951-:8],1'b0})+$signed(-{in[959-:8],2'b0})+$signed(sharing14)+$signed(1);
assign weighted_sum[186] = $signed({in[967-:8],1'b0})+$signed(-{in[975-:8],2'b0})+$signed(-{in[983-:8],2'b0})+$signed(-in[535-:8])+$signed({in[743-:8],1'b0})+$signed(in[743-:8])+$signed(-{in[759-:8],2'b0})+$signed(sharing15)+$signed(1);
assign weighted_sum[187] = $signed(-{in[775-:8],2'b0})+$signed({in[983-:8],1'b0})+$signed(-{in[991-:8],2'b0})+$signed(-{in[999-:8],2'b0})+$signed(-in[551-:8])+$signed({in[759-:8],1'b0})+$signed(in[759-:8])+$signed(sharing16)+$signed(1);
assign weighted_sum[188] = $signed({in[775-:8],1'b0})+$signed(in[775-:8])+$signed(-{in[791-:8],2'b0})+$signed({in[999-:8],1'b0})+$signed(-{in[1007-:8],2'b0})+$signed(-{in[1015-:8],2'b0})+$signed(-in[567-:8])+$signed(sharing17)+$signed(1);
assign weighted_sum[189] = $signed(-{in[1031-:8],2'b0})+$signed(-in[583-:8])+$signed({in[791-:8],1'b0})+$signed(in[791-:8])+$signed(-{in[807-:8],2'b0})+$signed({in[1015-:8],1'b0})+$signed(-{in[1023-:8],2'b0})+$signed(sharing18)+$signed(1);
assign weighted_sum[190] = $signed({in[1031-:8],1'b0})+$signed(-{in[1039-:8],2'b0})+$signed(-{in[1047-:8],2'b0})+$signed(-in[599-:8])+$signed({in[807-:8],1'b0})+$signed(in[807-:8])+$signed(-{in[823-:8],2'b0})+$signed(sharing19)+$signed(1);
assign weighted_sum[191] = $signed(-{in[839-:8],2'b0})+$signed({in[1047-:8],1'b0})+$signed(-{in[1055-:8],2'b0})+$signed(-{in[1063-:8],2'b0})+$signed(-in[615-:8])+$signed({in[823-:8],1'b0})+$signed(in[823-:8])+$signed(sharing150)+$signed(1);
assign weighted_sum[192] = $signed({in[839-:8],1'b0})+$signed(in[839-:8])+$signed(-{in[855-:8],2'b0})+$signed({in[1063-:8],1'b0})+$signed(-{in[1071-:8],2'b0})+$signed(-{in[1079-:8],2'b0})+$signed(-in[631-:8])+$signed(sharing20)+$signed(1);
assign weighted_sum[193] = $signed(-{in[1095-:8],2'b0})+$signed(-in[647-:8])+$signed({in[855-:8],1'b0})+$signed(in[855-:8])+$signed(-{in[871-:8],2'b0})+$signed({in[1079-:8],1'b0})+$signed(-{in[1087-:8],2'b0})+$signed(sharing21)+$signed(1);
assign weighted_sum[194] = $signed({in[1095-:8],1'b0})+$signed(-{in[1103-:8],2'b0})+$signed(-{in[1111-:8],2'b0})+$signed(-in[663-:8])+$signed({in[871-:8],1'b0})+$signed(in[871-:8])+$signed(-{in[887-:8],2'b0})+$signed(sharing22)+$signed(1);
assign weighted_sum[195] = $signed({in[1351-:8],1'b0})+$signed(-{in[1359-:8],2'b0})+$signed(-{in[1367-:8],2'b0})+$signed(-in[919-:8])+$signed({in[1127-:8],1'b0})+$signed(in[1127-:8])+$signed(-{in[1143-:8],2'b0})+$signed(sharing23)+$signed(1);
assign weighted_sum[196] = $signed(-{in[1159-:8],2'b0})+$signed({in[1367-:8],1'b0})+$signed(-{in[1375-:8],2'b0})+$signed(-{in[1383-:8],2'b0})+$signed(-in[935-:8])+$signed({in[1143-:8],1'b0})+$signed(in[1143-:8])+$signed(sharing24)+$signed(1);
assign weighted_sum[197] = $signed({in[1159-:8],1'b0})+$signed(in[1159-:8])+$signed(-{in[1175-:8],2'b0})+$signed({in[1383-:8],1'b0})+$signed(-{in[1391-:8],2'b0})+$signed(-{in[1399-:8],2'b0})+$signed(-in[951-:8])+$signed(sharing25)+$signed(1);
assign weighted_sum[198] = $signed(-{in[1415-:8],2'b0})+$signed(-in[967-:8])+$signed({in[1175-:8],1'b0})+$signed(in[1175-:8])+$signed(-{in[1191-:8],2'b0})+$signed({in[1399-:8],1'b0})+$signed(-{in[1407-:8],2'b0})+$signed(sharing26)+$signed(1);
assign weighted_sum[199] = $signed({in[1415-:8],1'b0})+$signed(-{in[1423-:8],2'b0})+$signed(-{in[1431-:8],2'b0})+$signed(-in[983-:8])+$signed({in[1191-:8],1'b0})+$signed(in[1191-:8])+$signed(-{in[1207-:8],2'b0})+$signed(sharing151)+$signed(1);
assign weighted_sum[200] = $signed(-{in[1223-:8],2'b0})+$signed({in[1431-:8],1'b0})+$signed(-{in[1439-:8],2'b0})+$signed(-{in[1447-:8],2'b0})+$signed(-in[999-:8])+$signed({in[1207-:8],1'b0})+$signed(in[1207-:8])+$signed(sharing27)+$signed(1);
assign weighted_sum[201] = $signed({in[1223-:8],1'b0})+$signed(in[1223-:8])+$signed(-{in[1239-:8],2'b0})+$signed({in[1447-:8],1'b0})+$signed(-{in[1455-:8],2'b0})+$signed(-{in[1463-:8],2'b0})+$signed(-in[1015-:8])+$signed(sharing28)+$signed(1);
assign weighted_sum[202] = $signed(-{in[1479-:8],2'b0})+$signed(-in[1031-:8])+$signed({in[1239-:8],1'b0})+$signed(in[1239-:8])+$signed(-{in[1255-:8],2'b0})+$signed({in[1463-:8],1'b0})+$signed(-{in[1471-:8],2'b0})+$signed(sharing29)+$signed(1);
assign weighted_sum[203] = $signed({in[1479-:8],1'b0})+$signed(-{in[1487-:8],2'b0})+$signed(-{in[1495-:8],2'b0})+$signed(-in[1047-:8])+$signed({in[1255-:8],1'b0})+$signed(in[1255-:8])+$signed(-{in[1271-:8],2'b0})+$signed(sharing30)+$signed(1);
assign weighted_sum[204] = $signed(-{in[1287-:8],2'b0})+$signed({in[1495-:8],1'b0})+$signed(-{in[1503-:8],2'b0})+$signed(-{in[1511-:8],2'b0})+$signed(-in[1063-:8])+$signed({in[1271-:8],1'b0})+$signed(in[1271-:8])+$signed(sharing31)+$signed(1);
assign weighted_sum[205] = $signed({in[1287-:8],1'b0})+$signed(in[1287-:8])+$signed(-{in[1303-:8],2'b0})+$signed({in[1511-:8],1'b0})+$signed(-{in[1519-:8],2'b0})+$signed(-{in[1527-:8],2'b0})+$signed(-in[1079-:8])+$signed(sharing32)+$signed(1);
assign weighted_sum[206] = $signed(-{in[1543-:8],2'b0})+$signed(-in[1095-:8])+$signed({in[1303-:8],1'b0})+$signed(in[1303-:8])+$signed(-{in[1319-:8],2'b0})+$signed({in[1527-:8],1'b0})+$signed(-{in[1535-:8],2'b0})+$signed(sharing33)+$signed(1);
assign weighted_sum[207] = $signed({in[1543-:8],1'b0})+$signed(-{in[1551-:8],2'b0})+$signed(-{in[1559-:8],2'b0})+$signed(-in[1111-:8])+$signed({in[1319-:8],1'b0})+$signed(in[1319-:8])+$signed(-{in[1335-:8],2'b0})+$signed(sharing152)+$signed(1);
assign weighted_sum[208] = $signed({in[1799-:8],1'b0})+$signed(-{in[1807-:8],2'b0})+$signed(-{in[1815-:8],2'b0})+$signed(-in[1367-:8])+$signed({in[1575-:8],1'b0})+$signed(in[1575-:8])+$signed(-{in[1591-:8],2'b0})+$signed(sharing34)+$signed(1);
assign weighted_sum[209] = $signed(-{in[1607-:8],2'b0})+$signed({in[1815-:8],1'b0})+$signed(-{in[1823-:8],2'b0})+$signed(-{in[1831-:8],2'b0})+$signed(-in[1383-:8])+$signed({in[1591-:8],1'b0})+$signed(in[1591-:8])+$signed(sharing35)+$signed(1);
assign weighted_sum[210] = $signed({in[1607-:8],1'b0})+$signed(in[1607-:8])+$signed(-{in[1623-:8],2'b0})+$signed({in[1831-:8],1'b0})+$signed(-{in[1839-:8],2'b0})+$signed(-{in[1847-:8],2'b0})+$signed(-in[1399-:8])+$signed(sharing36)+$signed(1);
assign weighted_sum[211] = $signed(-{in[1863-:8],2'b0})+$signed(-in[1415-:8])+$signed({in[1623-:8],1'b0})+$signed(in[1623-:8])+$signed(-{in[1639-:8],2'b0})+$signed({in[1847-:8],1'b0})+$signed(-{in[1855-:8],2'b0})+$signed(sharing37)+$signed(1);
assign weighted_sum[212] = $signed({in[1863-:8],1'b0})+$signed(-{in[1871-:8],2'b0})+$signed(-{in[1879-:8],2'b0})+$signed(-in[1431-:8])+$signed({in[1639-:8],1'b0})+$signed(in[1639-:8])+$signed(-{in[1655-:8],2'b0})+$signed(sharing38)+$signed(1);
assign weighted_sum[213] = $signed(-{in[1671-:8],2'b0})+$signed({in[1879-:8],1'b0})+$signed(-{in[1887-:8],2'b0})+$signed(-{in[1895-:8],2'b0})+$signed(-in[1447-:8])+$signed({in[1655-:8],1'b0})+$signed(in[1655-:8])+$signed(sharing39)+$signed(1);
assign weighted_sum[214] = $signed({in[1671-:8],1'b0})+$signed(in[1671-:8])+$signed(-{in[1687-:8],2'b0})+$signed({in[1895-:8],1'b0})+$signed(-{in[1903-:8],2'b0})+$signed(-{in[1911-:8],2'b0})+$signed(-in[1463-:8])+$signed(sharing40)+$signed(1);
assign weighted_sum[215] = $signed(-{in[1927-:8],2'b0})+$signed(-in[1479-:8])+$signed({in[1687-:8],1'b0})+$signed(in[1687-:8])+$signed(-{in[1703-:8],2'b0})+$signed({in[1911-:8],1'b0})+$signed(-{in[1919-:8],2'b0})+$signed(sharing153)+$signed(1);
assign weighted_sum[216] = $signed({in[1927-:8],1'b0})+$signed(-{in[1935-:8],2'b0})+$signed(-{in[1943-:8],2'b0})+$signed(-in[1495-:8])+$signed({in[1703-:8],1'b0})+$signed(in[1703-:8])+$signed(-{in[1719-:8],2'b0})+$signed(sharing41)+$signed(1);
assign weighted_sum[217] = $signed(-{in[1735-:8],2'b0})+$signed({in[1943-:8],1'b0})+$signed(-{in[1951-:8],2'b0})+$signed(-{in[1959-:8],2'b0})+$signed(-in[1511-:8])+$signed({in[1719-:8],1'b0})+$signed(in[1719-:8])+$signed(sharing42)+$signed(1);
assign weighted_sum[218] = $signed({in[1735-:8],1'b0})+$signed(in[1735-:8])+$signed(-{in[1751-:8],2'b0})+$signed({in[1959-:8],1'b0})+$signed(-{in[1967-:8],2'b0})+$signed(-{in[1975-:8],2'b0})+$signed(-in[1527-:8])+$signed(sharing43)+$signed(1);
assign weighted_sum[219] = $signed(-{in[1991-:8],2'b0})+$signed(-in[1543-:8])+$signed({in[1751-:8],1'b0})+$signed(in[1751-:8])+$signed(-{in[1767-:8],2'b0})+$signed({in[1975-:8],1'b0})+$signed(-{in[1983-:8],2'b0})+$signed(sharing44)+$signed(1);
assign weighted_sum[220] = $signed({in[1991-:8],1'b0})+$signed(-{in[1999-:8],2'b0})+$signed(-{in[2007-:8],2'b0})+$signed(-in[1559-:8])+$signed({in[1767-:8],1'b0})+$signed(in[1767-:8])+$signed(-{in[1783-:8],2'b0})+$signed(sharing45)+$signed(1);
assign weighted_sum[221] = $signed({in[2247-:8],1'b0})+$signed(-{in[2255-:8],2'b0})+$signed(-{in[2263-:8],2'b0})+$signed(-in[1815-:8])+$signed({in[2023-:8],1'b0})+$signed(in[2023-:8])+$signed(-{in[2039-:8],2'b0})+$signed(sharing46)+$signed(1);
assign weighted_sum[222] = $signed(-{in[2055-:8],2'b0})+$signed({in[2263-:8],1'b0})+$signed(-{in[2271-:8],2'b0})+$signed(-{in[2279-:8],2'b0})+$signed(-in[1831-:8])+$signed({in[2039-:8],1'b0})+$signed(in[2039-:8])+$signed(sharing47)+$signed(1);
assign weighted_sum[223] = $signed({in[2055-:8],1'b0})+$signed(in[2055-:8])+$signed(-{in[2071-:8],2'b0})+$signed({in[2279-:8],1'b0})+$signed(-{in[2287-:8],2'b0})+$signed(-{in[2295-:8],2'b0})+$signed(-in[1847-:8])+$signed(sharing154)+$signed(1);
assign weighted_sum[224] = $signed(-{in[2311-:8],2'b0})+$signed(-in[1863-:8])+$signed({in[2071-:8],1'b0})+$signed(in[2071-:8])+$signed(-{in[2087-:8],2'b0})+$signed({in[2295-:8],1'b0})+$signed(-{in[2303-:8],2'b0})+$signed(sharing48)+$signed(1);
assign weighted_sum[225] = $signed({in[2311-:8],1'b0})+$signed(-{in[2319-:8],2'b0})+$signed(-{in[2327-:8],2'b0})+$signed(-in[1879-:8])+$signed({in[2087-:8],1'b0})+$signed(in[2087-:8])+$signed(-{in[2103-:8],2'b0})+$signed(sharing49)+$signed(1);
assign weighted_sum[226] = $signed(-{in[2119-:8],2'b0})+$signed({in[2327-:8],1'b0})+$signed(-{in[2335-:8],2'b0})+$signed(-{in[2343-:8],2'b0})+$signed(-in[1895-:8])+$signed({in[2103-:8],1'b0})+$signed(in[2103-:8])+$signed(sharing50)+$signed(1);
assign weighted_sum[227] = $signed({in[2119-:8],1'b0})+$signed(in[2119-:8])+$signed(-{in[2135-:8],2'b0})+$signed({in[2343-:8],1'b0})+$signed(-{in[2351-:8],2'b0})+$signed(-{in[2359-:8],2'b0})+$signed(-in[1911-:8])+$signed(sharing51)+$signed(1);
assign weighted_sum[228] = $signed(-{in[2375-:8],2'b0})+$signed(-in[1927-:8])+$signed({in[2135-:8],1'b0})+$signed(in[2135-:8])+$signed(-{in[2151-:8],2'b0})+$signed({in[2359-:8],1'b0})+$signed(-{in[2367-:8],2'b0})+$signed(sharing52)+$signed(1);
assign weighted_sum[229] = $signed({in[2375-:8],1'b0})+$signed(-{in[2383-:8],2'b0})+$signed(-{in[2391-:8],2'b0})+$signed(-in[1943-:8])+$signed({in[2151-:8],1'b0})+$signed(in[2151-:8])+$signed(-{in[2167-:8],2'b0})+$signed(sharing53)+$signed(1);
assign weighted_sum[230] = $signed(-{in[2183-:8],2'b0})+$signed({in[2391-:8],1'b0})+$signed(-{in[2399-:8],2'b0})+$signed(-{in[2407-:8],2'b0})+$signed(-in[1959-:8])+$signed({in[2167-:8],1'b0})+$signed(in[2167-:8])+$signed(sharing54)+$signed(1);
assign weighted_sum[231] = $signed({in[2183-:8],1'b0})+$signed(in[2183-:8])+$signed(-{in[2199-:8],2'b0})+$signed({in[2407-:8],1'b0})+$signed(-{in[2415-:8],2'b0})+$signed(-{in[2423-:8],2'b0})+$signed(-in[1975-:8])+$signed(sharing155)+$signed(1);
assign weighted_sum[232] = $signed(-{in[2439-:8],2'b0})+$signed(-in[1991-:8])+$signed({in[2199-:8],1'b0})+$signed(in[2199-:8])+$signed(-{in[2215-:8],2'b0})+$signed({in[2423-:8],1'b0})+$signed(-{in[2431-:8],2'b0})+$signed(sharing55)+$signed(1);
assign weighted_sum[233] = $signed({in[2439-:8],1'b0})+$signed(-{in[2447-:8],2'b0})+$signed(-{in[2455-:8],2'b0})+$signed(-in[2007-:8])+$signed({in[2215-:8],1'b0})+$signed(in[2215-:8])+$signed(-{in[2231-:8],2'b0})+$signed(sharing56)+$signed(1);
assign weighted_sum[234] = $signed({in[2695-:8],1'b0})+$signed(-{in[2703-:8],2'b0})+$signed(-{in[2711-:8],2'b0})+$signed(-in[2263-:8])+$signed({in[2471-:8],1'b0})+$signed(in[2471-:8])+$signed(-{in[2487-:8],2'b0})+$signed(sharing57)+$signed(1);
assign weighted_sum[235] = $signed(-{in[2503-:8],2'b0})+$signed({in[2711-:8],1'b0})+$signed(-{in[2719-:8],2'b0})+$signed(-{in[2727-:8],2'b0})+$signed(-in[2279-:8])+$signed({in[2487-:8],1'b0})+$signed(in[2487-:8])+$signed(sharing58)+$signed(1);
assign weighted_sum[236] = $signed({in[2503-:8],1'b0})+$signed(in[2503-:8])+$signed(-{in[2519-:8],2'b0})+$signed({in[2727-:8],1'b0})+$signed(-{in[2735-:8],2'b0})+$signed(-{in[2743-:8],2'b0})+$signed(-in[2295-:8])+$signed(sharing59)+$signed(1);
assign weighted_sum[237] = $signed(-{in[2759-:8],2'b0})+$signed(-in[2311-:8])+$signed({in[2519-:8],1'b0})+$signed(in[2519-:8])+$signed(-{in[2535-:8],2'b0})+$signed({in[2743-:8],1'b0})+$signed(-{in[2751-:8],2'b0})+$signed(sharing60)+$signed(1);
assign weighted_sum[238] = $signed({in[2759-:8],1'b0})+$signed(-{in[2767-:8],2'b0})+$signed(-{in[2775-:8],2'b0})+$signed(-in[2327-:8])+$signed({in[2535-:8],1'b0})+$signed(in[2535-:8])+$signed(-{in[2551-:8],2'b0})+$signed(sharing61)+$signed(1);
assign weighted_sum[239] = $signed(-{in[2567-:8],2'b0})+$signed({in[2775-:8],1'b0})+$signed(-{in[2783-:8],2'b0})+$signed(-{in[2791-:8],2'b0})+$signed(-in[2343-:8])+$signed({in[2551-:8],1'b0})+$signed(in[2551-:8])+$signed(sharing156)+$signed(1);
assign weighted_sum[240] = $signed({in[2567-:8],1'b0})+$signed(in[2567-:8])+$signed(-{in[2583-:8],2'b0})+$signed({in[2791-:8],1'b0})+$signed(-{in[2799-:8],2'b0})+$signed(-{in[2807-:8],2'b0})+$signed(-in[2359-:8])+$signed(sharing62)+$signed(1);
assign weighted_sum[241] = $signed(-{in[2823-:8],2'b0})+$signed(-in[2375-:8])+$signed({in[2583-:8],1'b0})+$signed(in[2583-:8])+$signed(-{in[2599-:8],2'b0})+$signed({in[2807-:8],1'b0})+$signed(-{in[2815-:8],2'b0})+$signed(sharing63)+$signed(1);
assign weighted_sum[242] = $signed({in[2823-:8],1'b0})+$signed(-{in[2831-:8],2'b0})+$signed(-{in[2839-:8],2'b0})+$signed(-in[2391-:8])+$signed({in[2599-:8],1'b0})+$signed(in[2599-:8])+$signed(-{in[2615-:8],2'b0})+$signed(sharing64)+$signed(1);
assign weighted_sum[243] = $signed(-{in[2631-:8],2'b0})+$signed({in[2839-:8],1'b0})+$signed(-{in[2847-:8],2'b0})+$signed(-{in[2855-:8],2'b0})+$signed(-in[2407-:8])+$signed({in[2615-:8],1'b0})+$signed(in[2615-:8])+$signed(sharing65)+$signed(1);
assign weighted_sum[244] = $signed({in[2631-:8],1'b0})+$signed(in[2631-:8])+$signed(-{in[2647-:8],2'b0})+$signed({in[2855-:8],1'b0})+$signed(-{in[2863-:8],2'b0})+$signed(-{in[2871-:8],2'b0})+$signed(-in[2423-:8])+$signed(sharing66)+$signed(1);
assign weighted_sum[245] = $signed(-{in[2887-:8],2'b0})+$signed(-in[2439-:8])+$signed({in[2647-:8],1'b0})+$signed(in[2647-:8])+$signed(-{in[2663-:8],2'b0})+$signed({in[2871-:8],1'b0})+$signed(-{in[2879-:8],2'b0})+$signed(sharing67)+$signed(1);
assign weighted_sum[246] = $signed({in[2887-:8],1'b0})+$signed(-{in[2895-:8],2'b0})+$signed(-{in[2903-:8],2'b0})+$signed(-in[2455-:8])+$signed({in[2663-:8],1'b0})+$signed(in[2663-:8])+$signed(-{in[2679-:8],2'b0})+$signed(sharing68)+$signed(1);
assign weighted_sum[247] = $signed({in[3143-:8],1'b0})+$signed(-{in[3151-:8],2'b0})+$signed(-{in[3159-:8],2'b0})+$signed(-in[2711-:8])+$signed({in[2919-:8],1'b0})+$signed(in[2919-:8])+$signed(-{in[2935-:8],2'b0})+$signed(sharing157)+$signed(1);
assign weighted_sum[248] = $signed(-{in[2951-:8],2'b0})+$signed({in[3159-:8],1'b0})+$signed(-{in[3167-:8],2'b0})+$signed(-{in[3175-:8],2'b0})+$signed(-in[2727-:8])+$signed({in[2935-:8],1'b0})+$signed(in[2935-:8])+$signed(sharing69)+$signed(1);
assign weighted_sum[249] = $signed({in[2951-:8],1'b0})+$signed(in[2951-:8])+$signed(-{in[2967-:8],2'b0})+$signed({in[3175-:8],1'b0})+$signed(-{in[3183-:8],2'b0})+$signed(-{in[3191-:8],2'b0})+$signed(-in[2743-:8])+$signed(sharing70)+$signed(1);
assign weighted_sum[250] = $signed(-{in[3207-:8],2'b0})+$signed(-in[2759-:8])+$signed({in[2967-:8],1'b0})+$signed(in[2967-:8])+$signed(-{in[2983-:8],2'b0})+$signed({in[3191-:8],1'b0})+$signed(-{in[3199-:8],2'b0})+$signed(sharing71)+$signed(1);
assign weighted_sum[251] = $signed({in[3207-:8],1'b0})+$signed(-{in[3215-:8],2'b0})+$signed(-{in[3223-:8],2'b0})+$signed(-in[2775-:8])+$signed({in[2983-:8],1'b0})+$signed(in[2983-:8])+$signed(-{in[2999-:8],2'b0})+$signed(sharing72)+$signed(1);
assign weighted_sum[252] = $signed(-{in[3015-:8],2'b0})+$signed({in[3223-:8],1'b0})+$signed(-{in[3231-:8],2'b0})+$signed(-{in[3239-:8],2'b0})+$signed(-in[2791-:8])+$signed({in[2999-:8],1'b0})+$signed(in[2999-:8])+$signed(sharing73)+$signed(1);
assign weighted_sum[253] = $signed({in[3015-:8],1'b0})+$signed(in[3015-:8])+$signed(-{in[3031-:8],2'b0})+$signed({in[3239-:8],1'b0})+$signed(-{in[3247-:8],2'b0})+$signed(-{in[3255-:8],2'b0})+$signed(-in[2807-:8])+$signed(sharing74)+$signed(1);
assign weighted_sum[254] = $signed(-{in[3271-:8],2'b0})+$signed(-in[2823-:8])+$signed({in[3031-:8],1'b0})+$signed(in[3031-:8])+$signed(-{in[3047-:8],2'b0})+$signed({in[3255-:8],1'b0})+$signed(-{in[3263-:8],2'b0})+$signed(sharing75)+$signed(1);
assign weighted_sum[255] = $signed({in[3271-:8],1'b0})+$signed(-{in[3279-:8],2'b0})+$signed(-{in[3287-:8],2'b0})+$signed(-in[2839-:8])+$signed({in[3047-:8],1'b0})+$signed(in[3047-:8])+$signed(-{in[3063-:8],2'b0})+$signed(sharing158)+$signed(1);
assign weighted_sum[256] = $signed(-{in[3079-:8],2'b0})+$signed({in[3287-:8],1'b0})+$signed(-{in[3295-:8],2'b0})+$signed(-{in[3303-:8],2'b0})+$signed(-in[2855-:8])+$signed({in[3063-:8],1'b0})+$signed(in[3063-:8])+$signed(sharing76)+$signed(1);
assign weighted_sum[257] = $signed({in[3079-:8],1'b0})+$signed(in[3079-:8])+$signed(-{in[3095-:8],2'b0})+$signed({in[3303-:8],1'b0})+$signed(-{in[3311-:8],2'b0})+$signed(-{in[3319-:8],2'b0})+$signed(-in[2871-:8])+$signed(sharing77)+$signed(1);
assign weighted_sum[258] = $signed(-{in[3335-:8],2'b0})+$signed(-in[2887-:8])+$signed({in[3095-:8],1'b0})+$signed(in[3095-:8])+$signed(-{in[3111-:8],2'b0})+$signed({in[3319-:8],1'b0})+$signed(-{in[3327-:8],2'b0})+$signed(sharing78)+$signed(1);
assign weighted_sum[259] = $signed({in[3335-:8],1'b0})+$signed(-{in[3343-:8],2'b0})+$signed(-{in[3351-:8],2'b0})+$signed(-in[2903-:8])+$signed({in[3111-:8],1'b0})+$signed(in[3111-:8])+$signed(-{in[3127-:8],2'b0})+$signed(sharing79)+$signed(1);
assign weighted_sum[260] = $signed({in[3591-:8],1'b0})+$signed(-{in[3599-:8],2'b0})+$signed(-{in[3607-:8],2'b0})+$signed(-in[3159-:8])+$signed({in[3367-:8],1'b0})+$signed(in[3367-:8])+$signed(-{in[3383-:8],2'b0})+$signed(sharing80)+$signed(1);
assign weighted_sum[261] = $signed(-{in[3399-:8],2'b0})+$signed({in[3607-:8],1'b0})+$signed(-{in[3615-:8],2'b0})+$signed(-{in[3623-:8],2'b0})+$signed(-in[3175-:8])+$signed({in[3383-:8],1'b0})+$signed(in[3383-:8])+$signed(sharing81)+$signed(1);
assign weighted_sum[262] = $signed({in[3399-:8],1'b0})+$signed(in[3399-:8])+$signed(-{in[3415-:8],2'b0})+$signed({in[3623-:8],1'b0})+$signed(-{in[3631-:8],2'b0})+$signed(-{in[3639-:8],2'b0})+$signed(-in[3191-:8])+$signed(sharing82)+$signed(1);
assign weighted_sum[263] = $signed(-{in[3655-:8],2'b0})+$signed(-in[3207-:8])+$signed({in[3415-:8],1'b0})+$signed(in[3415-:8])+$signed(-{in[3431-:8],2'b0})+$signed({in[3639-:8],1'b0})+$signed(-{in[3647-:8],2'b0})+$signed(sharing159)+$signed(1);
assign weighted_sum[264] = $signed({in[3655-:8],1'b0})+$signed(-{in[3663-:8],2'b0})+$signed(-{in[3671-:8],2'b0})+$signed(-in[3223-:8])+$signed({in[3431-:8],1'b0})+$signed(in[3431-:8])+$signed(-{in[3447-:8],2'b0})+$signed(sharing83)+$signed(1);
assign weighted_sum[265] = $signed(-{in[3463-:8],2'b0})+$signed({in[3671-:8],1'b0})+$signed(-{in[3679-:8],2'b0})+$signed(-{in[3687-:8],2'b0})+$signed(-in[3239-:8])+$signed({in[3447-:8],1'b0})+$signed(in[3447-:8])+$signed(sharing84)+$signed(1);
assign weighted_sum[266] = $signed({in[3463-:8],1'b0})+$signed(in[3463-:8])+$signed(-{in[3479-:8],2'b0})+$signed({in[3687-:8],1'b0})+$signed(-{in[3695-:8],2'b0})+$signed(-{in[3703-:8],2'b0})+$signed(-in[3255-:8])+$signed(sharing85)+$signed(1);
assign weighted_sum[267] = $signed(-{in[3719-:8],2'b0})+$signed(-in[3271-:8])+$signed({in[3479-:8],1'b0})+$signed(in[3479-:8])+$signed(-{in[3495-:8],2'b0})+$signed({in[3703-:8],1'b0})+$signed(-{in[3711-:8],2'b0})+$signed(sharing86)+$signed(1);
assign weighted_sum[268] = $signed({in[3719-:8],1'b0})+$signed(-{in[3727-:8],2'b0})+$signed(-{in[3735-:8],2'b0})+$signed(-in[3287-:8])+$signed({in[3495-:8],1'b0})+$signed(in[3495-:8])+$signed(-{in[3511-:8],2'b0})+$signed(sharing87)+$signed(1);
assign weighted_sum[269] = $signed(-{in[3527-:8],2'b0})+$signed({in[3735-:8],1'b0})+$signed(-{in[3743-:8],2'b0})+$signed(-{in[3751-:8],2'b0})+$signed(-in[3303-:8])+$signed({in[3511-:8],1'b0})+$signed(in[3511-:8])+$signed(sharing88)+$signed(1);
assign weighted_sum[270] = $signed({in[3527-:8],1'b0})+$signed(in[3527-:8])+$signed(-{in[3543-:8],2'b0})+$signed({in[3751-:8],1'b0})+$signed(-{in[3759-:8],2'b0})+$signed(-{in[3767-:8],2'b0})+$signed(-in[3319-:8])+$signed(sharing89)+$signed(1);
assign weighted_sum[271] = $signed(-{in[3783-:8],2'b0})+$signed(-in[3335-:8])+$signed({in[3543-:8],1'b0})+$signed(in[3543-:8])+$signed(-{in[3559-:8],2'b0})+$signed({in[3767-:8],1'b0})+$signed(-{in[3775-:8],2'b0})+$signed(sharing160)+$signed(1);
assign weighted_sum[272] = $signed({in[3783-:8],1'b0})+$signed(-{in[3791-:8],2'b0})+$signed(-{in[3799-:8],2'b0})+$signed(-in[3351-:8])+$signed({in[3559-:8],1'b0})+$signed(in[3559-:8])+$signed(-{in[3575-:8],2'b0})+$signed(sharing90)+$signed(1);
assign weighted_sum[273] = $signed({in[4039-:8],1'b0})+$signed(-{in[4047-:8],2'b0})+$signed(-{in[4055-:8],2'b0})+$signed(-in[3607-:8])+$signed({in[3815-:8],1'b0})+$signed(in[3815-:8])+$signed(-{in[3831-:8],2'b0})+$signed(sharing91)+$signed(1);
assign weighted_sum[274] = $signed(-{in[3847-:8],2'b0})+$signed({in[4055-:8],1'b0})+$signed(-{in[4063-:8],2'b0})+$signed(-{in[4071-:8],2'b0})+$signed(-in[3623-:8])+$signed({in[3831-:8],1'b0})+$signed(in[3831-:8])+$signed(sharing92)+$signed(1);
assign weighted_sum[275] = $signed({in[3847-:8],1'b0})+$signed(in[3847-:8])+$signed(-{in[3863-:8],2'b0})+$signed({in[4071-:8],1'b0})+$signed(-{in[4079-:8],2'b0})+$signed(-{in[4087-:8],2'b0})+$signed(-in[3639-:8])+$signed(sharing93)+$signed(1);
assign weighted_sum[276] = $signed(-{in[4103-:8],2'b0})+$signed(-in[3655-:8])+$signed({in[3863-:8],1'b0})+$signed(in[3863-:8])+$signed(-{in[3879-:8],2'b0})+$signed({in[4087-:8],1'b0})+$signed(-{in[4095-:8],2'b0})+$signed(sharing94)+$signed(1);
assign weighted_sum[277] = $signed({in[4103-:8],1'b0})+$signed(-{in[4111-:8],2'b0})+$signed(-{in[4119-:8],2'b0})+$signed(-in[3671-:8])+$signed({in[3879-:8],1'b0})+$signed(in[3879-:8])+$signed(-{in[3895-:8],2'b0})+$signed(sharing95)+$signed(1);
assign weighted_sum[278] = $signed(-{in[3911-:8],2'b0})+$signed({in[4119-:8],1'b0})+$signed(-{in[4127-:8],2'b0})+$signed(-{in[4135-:8],2'b0})+$signed(-in[3687-:8])+$signed({in[3895-:8],1'b0})+$signed(in[3895-:8])+$signed(sharing96)+$signed(1);
assign weighted_sum[279] = $signed({in[3911-:8],1'b0})+$signed(in[3911-:8])+$signed(-{in[3927-:8],2'b0})+$signed({in[4135-:8],1'b0})+$signed(-{in[4143-:8],2'b0})+$signed(-{in[4151-:8],2'b0})+$signed(-in[3703-:8])+$signed(sharing161)+$signed(1);
assign weighted_sum[280] = $signed(-{in[4167-:8],2'b0})+$signed(-in[3719-:8])+$signed({in[3927-:8],1'b0})+$signed(in[3927-:8])+$signed(-{in[3943-:8],2'b0})+$signed({in[4151-:8],1'b0})+$signed(-{in[4159-:8],2'b0})+$signed(sharing97)+$signed(1);
assign weighted_sum[281] = $signed({in[4167-:8],1'b0})+$signed(-{in[4175-:8],2'b0})+$signed(-{in[4183-:8],2'b0})+$signed(-in[3735-:8])+$signed({in[3943-:8],1'b0})+$signed(in[3943-:8])+$signed(-{in[3959-:8],2'b0})+$signed(sharing98)+$signed(1);
assign weighted_sum[282] = $signed(-{in[3975-:8],2'b0})+$signed({in[4183-:8],1'b0})+$signed(-{in[4191-:8],2'b0})+$signed(-{in[4199-:8],2'b0})+$signed(-in[3751-:8])+$signed({in[3959-:8],1'b0})+$signed(in[3959-:8])+$signed(sharing99)+$signed(1);
assign weighted_sum[283] = $signed({in[3975-:8],1'b0})+$signed(in[3975-:8])+$signed(-{in[3991-:8],2'b0})+$signed({in[4199-:8],1'b0})+$signed(-{in[4207-:8],2'b0})+$signed(-{in[4215-:8],2'b0})+$signed(-in[3767-:8])+$signed(sharing100)+$signed(1);
assign weighted_sum[284] = $signed(-{in[4231-:8],2'b0})+$signed(-in[3783-:8])+$signed({in[3991-:8],1'b0})+$signed(in[3991-:8])+$signed(-{in[4007-:8],2'b0})+$signed({in[4215-:8],1'b0})+$signed(-{in[4223-:8],2'b0})+$signed(sharing101)+$signed(1);
assign weighted_sum[285] = $signed({in[4231-:8],1'b0})+$signed(-{in[4239-:8],2'b0})+$signed(-{in[4247-:8],2'b0})+$signed(-in[3799-:8])+$signed({in[4007-:8],1'b0})+$signed(in[4007-:8])+$signed(-{in[4023-:8],2'b0})+$signed(sharing102)+$signed(1);
assign weighted_sum[286] = $signed({in[4487-:8],1'b0})+$signed(-{in[4495-:8],2'b0})+$signed(-{in[4503-:8],2'b0})+$signed(-in[4055-:8])+$signed({in[4263-:8],1'b0})+$signed(in[4263-:8])+$signed(-{in[4279-:8],2'b0})+$signed(sharing103)+$signed(1);
assign weighted_sum[287] = $signed(-{in[4295-:8],2'b0})+$signed({in[4503-:8],1'b0})+$signed(-{in[4511-:8],2'b0})+$signed(-{in[4519-:8],2'b0})+$signed(-in[4071-:8])+$signed({in[4279-:8],1'b0})+$signed(in[4279-:8])+$signed(sharing162)+$signed(1);
assign weighted_sum[288] = $signed({in[4295-:8],1'b0})+$signed(in[4295-:8])+$signed(-{in[4311-:8],2'b0})+$signed({in[4519-:8],1'b0})+$signed(-{in[4527-:8],2'b0})+$signed(-{in[4535-:8],2'b0})+$signed(-in[4087-:8])+$signed(sharing104)+$signed(1);
assign weighted_sum[289] = $signed(-{in[4551-:8],2'b0})+$signed(-in[4103-:8])+$signed({in[4311-:8],1'b0})+$signed(in[4311-:8])+$signed(-{in[4327-:8],2'b0})+$signed({in[4535-:8],1'b0})+$signed(-{in[4543-:8],2'b0})+$signed(sharing105)+$signed(1);
assign weighted_sum[290] = $signed({in[4551-:8],1'b0})+$signed(-{in[4559-:8],2'b0})+$signed(-{in[4567-:8],2'b0})+$signed(-in[4119-:8])+$signed({in[4327-:8],1'b0})+$signed(in[4327-:8])+$signed(-{in[4343-:8],2'b0})+$signed(sharing106)+$signed(1);
assign weighted_sum[291] = $signed(-{in[4359-:8],2'b0})+$signed({in[4567-:8],1'b0})+$signed(-{in[4575-:8],2'b0})+$signed(-{in[4583-:8],2'b0})+$signed(-in[4135-:8])+$signed({in[4343-:8],1'b0})+$signed(in[4343-:8])+$signed(sharing107)+$signed(1);
assign weighted_sum[292] = $signed({in[4359-:8],1'b0})+$signed(in[4359-:8])+$signed(-{in[4375-:8],2'b0})+$signed({in[4583-:8],1'b0})+$signed(-{in[4591-:8],2'b0})+$signed(-{in[4599-:8],2'b0})+$signed(-in[4151-:8])+$signed(sharing108)+$signed(1);
assign weighted_sum[293] = $signed(-{in[4615-:8],2'b0})+$signed(-in[4167-:8])+$signed({in[4375-:8],1'b0})+$signed(in[4375-:8])+$signed(-{in[4391-:8],2'b0})+$signed({in[4599-:8],1'b0})+$signed(-{in[4607-:8],2'b0})+$signed(sharing109)+$signed(1);
assign weighted_sum[294] = $signed({in[4615-:8],1'b0})+$signed(-{in[4623-:8],2'b0})+$signed(-{in[4631-:8],2'b0})+$signed(-in[4183-:8])+$signed({in[4391-:8],1'b0})+$signed(in[4391-:8])+$signed(-{in[4407-:8],2'b0})+$signed(sharing110)+$signed(1);
assign weighted_sum[295] = $signed(-{in[4423-:8],2'b0})+$signed({in[4631-:8],1'b0})+$signed(-{in[4639-:8],2'b0})+$signed(-{in[4647-:8],2'b0})+$signed(-in[4199-:8])+$signed({in[4407-:8],1'b0})+$signed(in[4407-:8])+$signed(sharing163)+$signed(1);
assign weighted_sum[296] = $signed({in[4423-:8],1'b0})+$signed(in[4423-:8])+$signed(-{in[4439-:8],2'b0})+$signed({in[4647-:8],1'b0})+$signed(-{in[4655-:8],2'b0})+$signed(-{in[4663-:8],2'b0})+$signed(-in[4215-:8])+$signed(sharing111)+$signed(1);
assign weighted_sum[297] = $signed(-{in[4679-:8],2'b0})+$signed(-in[4231-:8])+$signed({in[4439-:8],1'b0})+$signed(in[4439-:8])+$signed(-{in[4455-:8],2'b0})+$signed({in[4663-:8],1'b0})+$signed(-{in[4671-:8],2'b0})+$signed(sharing112)+$signed(1);
assign weighted_sum[298] = $signed({in[4679-:8],1'b0})+$signed(-{in[4687-:8],2'b0})+$signed(-{in[4695-:8],2'b0})+$signed(-in[4247-:8])+$signed({in[4455-:8],1'b0})+$signed(in[4455-:8])+$signed(-{in[4471-:8],2'b0})+$signed(sharing113)+$signed(1);
assign weighted_sum[299] = $signed({in[4935-:8],1'b0})+$signed(-{in[4943-:8],2'b0})+$signed(-{in[4951-:8],2'b0})+$signed(-in[4503-:8])+$signed({in[4711-:8],1'b0})+$signed(in[4711-:8])+$signed(-{in[4727-:8],2'b0})+$signed(sharing114)+$signed(1);
assign weighted_sum[300] = $signed(-{in[4743-:8],2'b0})+$signed({in[4951-:8],1'b0})+$signed(-{in[4959-:8],2'b0})+$signed(-{in[4967-:8],2'b0})+$signed(-in[4519-:8])+$signed({in[4727-:8],1'b0})+$signed(in[4727-:8])+$signed(sharing115)+$signed(1);
assign weighted_sum[301] = $signed({in[4743-:8],1'b0})+$signed(in[4743-:8])+$signed(-{in[4759-:8],2'b0})+$signed({in[4967-:8],1'b0})+$signed(-{in[4975-:8],2'b0})+$signed(-{in[4983-:8],2'b0})+$signed(-in[4535-:8])+$signed(sharing116)+$signed(1);
assign weighted_sum[302] = $signed(-{in[4999-:8],2'b0})+$signed(-in[4551-:8])+$signed({in[4759-:8],1'b0})+$signed(in[4759-:8])+$signed(-{in[4775-:8],2'b0})+$signed({in[4983-:8],1'b0})+$signed(-{in[4991-:8],2'b0})+$signed(sharing117)+$signed(1);
assign weighted_sum[303] = $signed({in[4999-:8],1'b0})+$signed(-{in[5007-:8],2'b0})+$signed(-{in[5015-:8],2'b0})+$signed(-in[4567-:8])+$signed({in[4775-:8],1'b0})+$signed(in[4775-:8])+$signed(-{in[4791-:8],2'b0})+$signed(sharing164)+$signed(1);
assign weighted_sum[304] = $signed(-{in[4807-:8],2'b0})+$signed({in[5015-:8],1'b0})+$signed(-{in[5023-:8],2'b0})+$signed(-{in[5031-:8],2'b0})+$signed(-in[4583-:8])+$signed({in[4791-:8],1'b0})+$signed(in[4791-:8])+$signed(sharing118)+$signed(1);
assign weighted_sum[305] = $signed({in[4807-:8],1'b0})+$signed(in[4807-:8])+$signed(-{in[4823-:8],2'b0})+$signed({in[5031-:8],1'b0})+$signed(-{in[5039-:8],2'b0})+$signed(-{in[5047-:8],2'b0})+$signed(-in[4599-:8])+$signed(sharing119)+$signed(1);
assign weighted_sum[306] = $signed(-{in[5063-:8],2'b0})+$signed(-in[4615-:8])+$signed({in[4823-:8],1'b0})+$signed(in[4823-:8])+$signed(-{in[4839-:8],2'b0})+$signed({in[5047-:8],1'b0})+$signed(-{in[5055-:8],2'b0})+$signed(sharing120)+$signed(1);
assign weighted_sum[307] = $signed({in[5063-:8],1'b0})+$signed(-{in[5071-:8],2'b0})+$signed(-{in[5079-:8],2'b0})+$signed(-in[4631-:8])+$signed({in[4839-:8],1'b0})+$signed(in[4839-:8])+$signed(-{in[4855-:8],2'b0})+$signed(sharing121)+$signed(1);
assign weighted_sum[308] = $signed(-{in[4871-:8],2'b0})+$signed({in[5079-:8],1'b0})+$signed(-{in[5087-:8],2'b0})+$signed(-{in[5095-:8],2'b0})+$signed(-in[4647-:8])+$signed({in[4855-:8],1'b0})+$signed(in[4855-:8])+$signed(sharing122)+$signed(1);
assign weighted_sum[309] = $signed({in[4871-:8],1'b0})+$signed(in[4871-:8])+$signed(-{in[4887-:8],2'b0})+$signed({in[5095-:8],1'b0})+$signed(-{in[5103-:8],2'b0})+$signed(-{in[5111-:8],2'b0})+$signed(-in[4663-:8])+$signed(sharing123)+$signed(1);
assign weighted_sum[310] = $signed(-{in[5127-:8],2'b0})+$signed(-in[4679-:8])+$signed({in[4887-:8],1'b0})+$signed(in[4887-:8])+$signed(-{in[4903-:8],2'b0})+$signed({in[5111-:8],1'b0})+$signed(-{in[5119-:8],2'b0})+$signed(sharing124)+$signed(1);
assign weighted_sum[311] = $signed({in[5127-:8],1'b0})+$signed(-{in[5135-:8],2'b0})+$signed(-{in[5143-:8],2'b0})+$signed(-in[4695-:8])+$signed({in[4903-:8],1'b0})+$signed(in[4903-:8])+$signed(-{in[4919-:8],2'b0})+$signed(sharing165)+$signed(1);
assign weighted_sum[312] = $signed({in[5383-:8],1'b0})+$signed(-{in[5391-:8],2'b0})+$signed(-{in[5399-:8],2'b0})+$signed(-in[4951-:8])+$signed({in[5159-:8],1'b0})+$signed(in[5159-:8])+$signed(-{in[5175-:8],2'b0})+$signed(sharing125)+$signed(1);
assign weighted_sum[313] = $signed(-{in[5191-:8],2'b0})+$signed({in[5399-:8],1'b0})+$signed(-{in[5407-:8],2'b0})+$signed(-{in[5415-:8],2'b0})+$signed(-in[4967-:8])+$signed({in[5175-:8],1'b0})+$signed(in[5175-:8])+$signed(sharing126)+$signed(1);
assign weighted_sum[314] = $signed({in[5191-:8],1'b0})+$signed(in[5191-:8])+$signed(-{in[5207-:8],2'b0})+$signed({in[5415-:8],1'b0})+$signed(-{in[5423-:8],2'b0})+$signed(-{in[5431-:8],2'b0})+$signed(-in[4983-:8])+$signed(sharing127)+$signed(1);
assign weighted_sum[315] = $signed(-{in[5447-:8],2'b0})+$signed(-in[4999-:8])+$signed({in[5207-:8],1'b0})+$signed(in[5207-:8])+$signed(-{in[5223-:8],2'b0})+$signed({in[5431-:8],1'b0})+$signed(-{in[5439-:8],2'b0})+$signed(sharing128)+$signed(1);
assign weighted_sum[316] = $signed({in[5447-:8],1'b0})+$signed(-{in[5455-:8],2'b0})+$signed(-{in[5463-:8],2'b0})+$signed(-in[5015-:8])+$signed({in[5223-:8],1'b0})+$signed(in[5223-:8])+$signed(-{in[5239-:8],2'b0})+$signed(sharing129)+$signed(1);
assign weighted_sum[317] = $signed(-{in[5255-:8],2'b0})+$signed({in[5463-:8],1'b0})+$signed(-{in[5471-:8],2'b0})+$signed(-{in[5479-:8],2'b0})+$signed(-in[5031-:8])+$signed({in[5239-:8],1'b0})+$signed(in[5239-:8])+$signed(sharing130)+$signed(1);
assign weighted_sum[318] = $signed({in[5255-:8],1'b0})+$signed(in[5255-:8])+$signed(-{in[5271-:8],2'b0})+$signed({in[5479-:8],1'b0})+$signed(-{in[5487-:8],2'b0})+$signed(-{in[5495-:8],2'b0})+$signed(-in[5047-:8])+$signed(sharing131)+$signed(1);
assign weighted_sum[319] = $signed(-{in[5511-:8],2'b0})+$signed(-in[5063-:8])+$signed({in[5271-:8],1'b0})+$signed(in[5271-:8])+$signed(-{in[5287-:8],2'b0})+$signed({in[5495-:8],1'b0})+$signed(-{in[5503-:8],2'b0})+$signed(sharing166)+$signed(1);
assign weighted_sum[320] = $signed({in[5511-:8],1'b0})+$signed(-{in[5519-:8],2'b0})+$signed(-{in[5527-:8],2'b0})+$signed(-in[5079-:8])+$signed({in[5287-:8],1'b0})+$signed(in[5287-:8])+$signed(-{in[5303-:8],2'b0})+$signed(sharing132)+$signed(1);
assign weighted_sum[321] = $signed(-{in[5319-:8],2'b0})+$signed({in[5527-:8],1'b0})+$signed(-{in[5535-:8],2'b0})+$signed(-{in[5543-:8],2'b0})+$signed(-in[5095-:8])+$signed({in[5303-:8],1'b0})+$signed(in[5303-:8])+$signed(sharing133)+$signed(1);
assign weighted_sum[322] = $signed({in[5319-:8],1'b0})+$signed(in[5319-:8])+$signed(-{in[5335-:8],2'b0})+$signed({in[5543-:8],1'b0})+$signed(-{in[5551-:8],2'b0})+$signed(-{in[5559-:8],2'b0})+$signed(-in[5111-:8])+$signed(sharing134)+$signed(1);
assign weighted_sum[323] = $signed(-{in[5575-:8],2'b0})+$signed(-in[5127-:8])+$signed({in[5335-:8],1'b0})+$signed(in[5335-:8])+$signed(-{in[5351-:8],2'b0})+$signed({in[5559-:8],1'b0})+$signed(-{in[5567-:8],2'b0})+$signed(sharing135)+$signed(1);
assign weighted_sum[324] = $signed({in[5575-:8],1'b0})+$signed(-{in[5583-:8],2'b0})+$signed(-{in[5591-:8],2'b0})+$signed(-in[5143-:8])+$signed({in[5351-:8],1'b0})+$signed(in[5351-:8])+$signed(-{in[5367-:8],2'b0})+$signed(sharing136)+$signed(1);
assign weighted_sum[325] = $signed({in[5831-:8],1'b0})+$signed(-{in[5839-:8],2'b0})+$signed(-{in[5847-:8],2'b0})+$signed(-in[5399-:8])+$signed({in[5607-:8],1'b0})+$signed(in[5607-:8])+$signed(-{in[5623-:8],2'b0})+$signed(sharing137)+$signed(1);
assign weighted_sum[326] = $signed(-{in[5639-:8],2'b0})+$signed({in[5847-:8],1'b0})+$signed(-{in[5855-:8],2'b0})+$signed(-{in[5863-:8],2'b0})+$signed(-in[5415-:8])+$signed({in[5623-:8],1'b0})+$signed(in[5623-:8])+$signed(sharing138)+$signed(1);
assign weighted_sum[327] = $signed({in[5639-:8],1'b0})+$signed(in[5639-:8])+$signed(-{in[5655-:8],2'b0})+$signed({in[5863-:8],1'b0})+$signed(-{in[5871-:8],2'b0})+$signed(-{in[5879-:8],2'b0})+$signed(-in[5431-:8])+$signed(sharing167)+$signed(1);
assign weighted_sum[328] = $signed(-{in[5895-:8],2'b0})+$signed(-in[5447-:8])+$signed({in[5655-:8],1'b0})+$signed(in[5655-:8])+$signed(-{in[5671-:8],2'b0})+$signed({in[5879-:8],1'b0})+$signed(-{in[5887-:8],2'b0})+$signed(sharing139)+$signed(1);
assign weighted_sum[329] = $signed({in[5895-:8],1'b0})+$signed(-{in[5903-:8],2'b0})+$signed(-{in[5911-:8],2'b0})+$signed(-in[5463-:8])+$signed({in[5671-:8],1'b0})+$signed(in[5671-:8])+$signed(-{in[5687-:8],2'b0})+$signed(sharing140)+$signed(1);
assign weighted_sum[330] = $signed(-{in[5703-:8],2'b0})+$signed({in[5911-:8],1'b0})+$signed(-{in[5919-:8],2'b0})+$signed(-{in[5927-:8],2'b0})+$signed(-in[5479-:8])+$signed({in[5687-:8],1'b0})+$signed(in[5687-:8])+$signed(sharing141)+$signed(1);
assign weighted_sum[331] = $signed({in[5703-:8],1'b0})+$signed(in[5703-:8])+$signed(-{in[5719-:8],2'b0})+$signed({in[5927-:8],1'b0})+$signed(-{in[5935-:8],2'b0})+$signed(-{in[5943-:8],2'b0})+$signed(-in[5495-:8])+$signed(sharing142)+$signed(1);
assign weighted_sum[332] = $signed(-{in[5959-:8],2'b0})+$signed(-in[5511-:8])+$signed({in[5719-:8],1'b0})+$signed(in[5719-:8])+$signed(-{in[5735-:8],2'b0})+$signed({in[5943-:8],1'b0})+$signed(-{in[5951-:8],2'b0})+$signed(sharing143)+$signed(1);
assign weighted_sum[333] = $signed({in[5959-:8],1'b0})+$signed(-{in[5967-:8],2'b0})+$signed(-{in[5975-:8],2'b0})+$signed(-in[5527-:8])+$signed({in[5735-:8],1'b0})+$signed(in[5735-:8])+$signed(-{in[5751-:8],2'b0})+$signed(sharing144)+$signed(1);
assign weighted_sum[334] = $signed(-{in[5767-:8],2'b0})+$signed({in[5975-:8],1'b0})+$signed(-{in[5983-:8],2'b0})+$signed(-{in[5991-:8],2'b0})+$signed(-in[5543-:8])+$signed({in[5751-:8],1'b0})+$signed(in[5751-:8])+$signed(sharing145)+$signed(1);
assign weighted_sum[335] = $signed({in[5767-:8],1'b0})+$signed(in[5767-:8])+$signed(-{in[5783-:8],2'b0})+$signed({in[5991-:8],1'b0})+$signed(-{in[5999-:8],2'b0})+$signed(-{in[6007-:8],2'b0})+$signed(-in[5559-:8])+$signed(sharing168)+$signed(1);
assign weighted_sum[336] = $signed(-{in[6023-:8],2'b0})+$signed(-in[5575-:8])+$signed({in[5783-:8],1'b0})+$signed(in[5783-:8])+$signed(-{in[5799-:8],2'b0})+$signed({in[6007-:8],1'b0})+$signed(-{in[6015-:8],2'b0})+$signed(sharing146)+$signed(1);
assign weighted_sum[337] = $signed({in[6023-:8],1'b0})+$signed(-{in[6031-:8],2'b0})+$signed(-{in[6039-:8],2'b0})+$signed(-in[5591-:8])+$signed({in[5799-:8],1'b0})+$signed(in[5799-:8])+$signed(-{in[5815-:8],2'b0})+$signed(sharing147)+$signed(1);
assign weighted_sum[338] = $signed(-{in[455-:8],3'b0})+$signed(-{in[463-:8],3'b0})+$signed({in[15-:8],1'b0})+$signed({in[23-:8],2'b0})+$signed(-{in[471-:8],1'b0})+$signed(in[23-:8])+$signed(-{in[231-:8],2'b0})+$signed({in[239-:8],1'b0})+$signed({in[247-:8],1'b0})+$signed(in[247-:8])+$signed(sharing0)+$signed(-1);
assign weighted_sum[339] = $signed({in[263-:8],1'b0})+$signed(in[263-:8])+$signed(-{in[471-:8],3'b0})+$signed(-{in[479-:8],3'b0})+$signed({in[31-:8],1'b0})+$signed({in[39-:8],2'b0})+$signed(-{in[487-:8],1'b0})+$signed(in[39-:8])+$signed(-{in[247-:8],2'b0})+$signed({in[255-:8],1'b0})+$signed(sharing1)+$signed(-1);
assign weighted_sum[340] = $signed(-{in[263-:8],2'b0})+$signed({in[271-:8],1'b0})+$signed({in[279-:8],1'b0})+$signed(in[279-:8])+$signed(-{in[487-:8],3'b0})+$signed(-{in[495-:8],3'b0})+$signed({in[47-:8],1'b0})+$signed({in[55-:8],2'b0})+$signed(-{in[503-:8],1'b0})+$signed(in[55-:8])+$signed(sharing2)+$signed(-1);
assign weighted_sum[341] = $signed({in[71-:8],2'b0})+$signed(-{in[519-:8],1'b0})+$signed(in[71-:8])+$signed(-{in[279-:8],2'b0})+$signed({in[287-:8],1'b0})+$signed({in[295-:8],1'b0})+$signed(in[295-:8])+$signed(-{in[503-:8],3'b0})+$signed(-{in[511-:8],3'b0})+$signed({in[63-:8],1'b0})+$signed(sharing3)+$signed(-1);
assign weighted_sum[342] = $signed(-{in[519-:8],3'b0})+$signed(-{in[527-:8],3'b0})+$signed({in[79-:8],1'b0})+$signed({in[87-:8],2'b0})+$signed(-{in[535-:8],1'b0})+$signed(in[87-:8])+$signed(-{in[295-:8],2'b0})+$signed({in[303-:8],1'b0})+$signed({in[311-:8],1'b0})+$signed(in[311-:8])+$signed(sharing4)+$signed(-1);
assign weighted_sum[343] = $signed({in[327-:8],1'b0})+$signed(in[327-:8])+$signed(-{in[535-:8],3'b0})+$signed(-{in[543-:8],3'b0})+$signed({in[95-:8],1'b0})+$signed({in[103-:8],2'b0})+$signed(-{in[551-:8],1'b0})+$signed(in[103-:8])+$signed(-{in[311-:8],2'b0})+$signed({in[319-:8],1'b0})+$signed(sharing5)+$signed(-1);
assign weighted_sum[344] = $signed(-{in[327-:8],2'b0})+$signed({in[335-:8],1'b0})+$signed({in[343-:8],1'b0})+$signed(in[343-:8])+$signed(-{in[551-:8],3'b0})+$signed(-{in[559-:8],3'b0})+$signed({in[111-:8],1'b0})+$signed({in[119-:8],2'b0})+$signed(-{in[567-:8],1'b0})+$signed(in[119-:8])+$signed(sharing148)+$signed(-1);
assign weighted_sum[345] = $signed({in[135-:8],2'b0})+$signed(-{in[583-:8],1'b0})+$signed(in[135-:8])+$signed(-{in[343-:8],2'b0})+$signed({in[351-:8],1'b0})+$signed({in[359-:8],1'b0})+$signed(in[359-:8])+$signed(-{in[567-:8],3'b0})+$signed(-{in[575-:8],3'b0})+$signed({in[127-:8],1'b0})+$signed(sharing6)+$signed(-1);
assign weighted_sum[346] = $signed(-{in[583-:8],3'b0})+$signed(-{in[591-:8],3'b0})+$signed({in[143-:8],1'b0})+$signed({in[151-:8],2'b0})+$signed(-{in[599-:8],1'b0})+$signed(in[151-:8])+$signed(-{in[359-:8],2'b0})+$signed({in[367-:8],1'b0})+$signed({in[375-:8],1'b0})+$signed(in[375-:8])+$signed(sharing7)+$signed(-1);
assign weighted_sum[347] = $signed({in[391-:8],1'b0})+$signed(in[391-:8])+$signed(-{in[599-:8],3'b0})+$signed(-{in[607-:8],3'b0})+$signed({in[159-:8],1'b0})+$signed({in[167-:8],2'b0})+$signed(-{in[615-:8],1'b0})+$signed(in[167-:8])+$signed(-{in[375-:8],2'b0})+$signed({in[383-:8],1'b0})+$signed(sharing8)+$signed(-1);
assign weighted_sum[348] = $signed(-{in[391-:8],2'b0})+$signed({in[399-:8],1'b0})+$signed({in[407-:8],1'b0})+$signed(in[407-:8])+$signed(-{in[615-:8],3'b0})+$signed(-{in[623-:8],3'b0})+$signed({in[175-:8],1'b0})+$signed({in[183-:8],2'b0})+$signed(-{in[631-:8],1'b0})+$signed(in[183-:8])+$signed(sharing9)+$signed(-1);
assign weighted_sum[349] = $signed({in[199-:8],2'b0})+$signed(-{in[647-:8],1'b0})+$signed(in[199-:8])+$signed(-{in[407-:8],2'b0})+$signed({in[415-:8],1'b0})+$signed({in[423-:8],1'b0})+$signed(in[423-:8])+$signed(-{in[631-:8],3'b0})+$signed(-{in[639-:8],3'b0})+$signed({in[191-:8],1'b0})+$signed(sharing10)+$signed(-1);
assign weighted_sum[350] = $signed(-{in[647-:8],3'b0})+$signed(-{in[655-:8],3'b0})+$signed({in[207-:8],1'b0})+$signed({in[215-:8],2'b0})+$signed(-{in[663-:8],1'b0})+$signed(in[215-:8])+$signed(-{in[423-:8],2'b0})+$signed({in[431-:8],1'b0})+$signed({in[439-:8],1'b0})+$signed(in[439-:8])+$signed(sharing11)+$signed(-1);
assign weighted_sum[351] = $signed(-{in[903-:8],3'b0})+$signed(-{in[911-:8],3'b0})+$signed({in[463-:8],1'b0})+$signed({in[471-:8],2'b0})+$signed(-{in[919-:8],1'b0})+$signed(in[471-:8])+$signed(-{in[679-:8],2'b0})+$signed({in[687-:8],1'b0})+$signed({in[695-:8],1'b0})+$signed(in[695-:8])+$signed(sharing12)+$signed(-1);
assign weighted_sum[352] = $signed({in[711-:8],1'b0})+$signed(in[711-:8])+$signed(-{in[919-:8],3'b0})+$signed(-{in[927-:8],3'b0})+$signed({in[479-:8],1'b0})+$signed({in[487-:8],2'b0})+$signed(-{in[935-:8],1'b0})+$signed(in[487-:8])+$signed(-{in[695-:8],2'b0})+$signed({in[703-:8],1'b0})+$signed(sharing149)+$signed(-1);
assign weighted_sum[353] = $signed(-{in[711-:8],2'b0})+$signed({in[719-:8],1'b0})+$signed({in[727-:8],1'b0})+$signed(in[727-:8])+$signed(-{in[935-:8],3'b0})+$signed(-{in[943-:8],3'b0})+$signed({in[495-:8],1'b0})+$signed({in[503-:8],2'b0})+$signed(-{in[951-:8],1'b0})+$signed(in[503-:8])+$signed(sharing13)+$signed(-1);
assign weighted_sum[354] = $signed({in[519-:8],2'b0})+$signed(-{in[967-:8],1'b0})+$signed(in[519-:8])+$signed(-{in[727-:8],2'b0})+$signed({in[735-:8],1'b0})+$signed({in[743-:8],1'b0})+$signed(in[743-:8])+$signed(-{in[951-:8],3'b0})+$signed(-{in[959-:8],3'b0})+$signed({in[511-:8],1'b0})+$signed(sharing14)+$signed(-1);
assign weighted_sum[355] = $signed(-{in[967-:8],3'b0})+$signed(-{in[975-:8],3'b0})+$signed({in[527-:8],1'b0})+$signed({in[535-:8],2'b0})+$signed(-{in[983-:8],1'b0})+$signed(in[535-:8])+$signed(-{in[743-:8],2'b0})+$signed({in[751-:8],1'b0})+$signed({in[759-:8],1'b0})+$signed(in[759-:8])+$signed(sharing15)+$signed(-1);
assign weighted_sum[356] = $signed({in[775-:8],1'b0})+$signed(in[775-:8])+$signed(-{in[983-:8],3'b0})+$signed(-{in[991-:8],3'b0})+$signed({in[543-:8],1'b0})+$signed({in[551-:8],2'b0})+$signed(-{in[999-:8],1'b0})+$signed(in[551-:8])+$signed(-{in[759-:8],2'b0})+$signed({in[767-:8],1'b0})+$signed(sharing16)+$signed(-1);
assign weighted_sum[357] = $signed(-{in[775-:8],2'b0})+$signed({in[783-:8],1'b0})+$signed({in[791-:8],1'b0})+$signed(in[791-:8])+$signed(-{in[999-:8],3'b0})+$signed(-{in[1007-:8],3'b0})+$signed({in[559-:8],1'b0})+$signed({in[567-:8],2'b0})+$signed(-{in[1015-:8],1'b0})+$signed(in[567-:8])+$signed(sharing17)+$signed(-1);
assign weighted_sum[358] = $signed({in[583-:8],2'b0})+$signed(-{in[1031-:8],1'b0})+$signed(in[583-:8])+$signed(-{in[791-:8],2'b0})+$signed({in[799-:8],1'b0})+$signed({in[807-:8],1'b0})+$signed(in[807-:8])+$signed(-{in[1015-:8],3'b0})+$signed(-{in[1023-:8],3'b0})+$signed({in[575-:8],1'b0})+$signed(sharing18)+$signed(-1);
assign weighted_sum[359] = $signed(-{in[1031-:8],3'b0})+$signed(-{in[1039-:8],3'b0})+$signed({in[591-:8],1'b0})+$signed({in[599-:8],2'b0})+$signed(-{in[1047-:8],1'b0})+$signed(in[599-:8])+$signed(-{in[807-:8],2'b0})+$signed({in[815-:8],1'b0})+$signed({in[823-:8],1'b0})+$signed(in[823-:8])+$signed(sharing19)+$signed(-1);
assign weighted_sum[360] = $signed({in[839-:8],1'b0})+$signed(in[839-:8])+$signed(-{in[1047-:8],3'b0})+$signed(-{in[1055-:8],3'b0})+$signed({in[607-:8],1'b0})+$signed({in[615-:8],2'b0})+$signed(-{in[1063-:8],1'b0})+$signed(in[615-:8])+$signed(-{in[823-:8],2'b0})+$signed({in[831-:8],1'b0})+$signed(sharing150)+$signed(-1);
assign weighted_sum[361] = $signed(-{in[839-:8],2'b0})+$signed({in[847-:8],1'b0})+$signed({in[855-:8],1'b0})+$signed(in[855-:8])+$signed(-{in[1063-:8],3'b0})+$signed(-{in[1071-:8],3'b0})+$signed({in[623-:8],1'b0})+$signed({in[631-:8],2'b0})+$signed(-{in[1079-:8],1'b0})+$signed(in[631-:8])+$signed(sharing20)+$signed(-1);
assign weighted_sum[362] = $signed({in[647-:8],2'b0})+$signed(-{in[1095-:8],1'b0})+$signed(in[647-:8])+$signed(-{in[855-:8],2'b0})+$signed({in[863-:8],1'b0})+$signed({in[871-:8],1'b0})+$signed(in[871-:8])+$signed(-{in[1079-:8],3'b0})+$signed(-{in[1087-:8],3'b0})+$signed({in[639-:8],1'b0})+$signed(sharing21)+$signed(-1);
assign weighted_sum[363] = $signed(-{in[1095-:8],3'b0})+$signed(-{in[1103-:8],3'b0})+$signed({in[655-:8],1'b0})+$signed({in[663-:8],2'b0})+$signed(-{in[1111-:8],1'b0})+$signed(in[663-:8])+$signed(-{in[871-:8],2'b0})+$signed({in[879-:8],1'b0})+$signed({in[887-:8],1'b0})+$signed(in[887-:8])+$signed(sharing22)+$signed(-1);
assign weighted_sum[364] = $signed(-{in[1351-:8],3'b0})+$signed(-{in[1359-:8],3'b0})+$signed({in[911-:8],1'b0})+$signed({in[919-:8],2'b0})+$signed(-{in[1367-:8],1'b0})+$signed(in[919-:8])+$signed(-{in[1127-:8],2'b0})+$signed({in[1135-:8],1'b0})+$signed({in[1143-:8],1'b0})+$signed(in[1143-:8])+$signed(sharing23)+$signed(-1);
assign weighted_sum[365] = $signed({in[1159-:8],1'b0})+$signed(in[1159-:8])+$signed(-{in[1367-:8],3'b0})+$signed(-{in[1375-:8],3'b0})+$signed({in[927-:8],1'b0})+$signed({in[935-:8],2'b0})+$signed(-{in[1383-:8],1'b0})+$signed(in[935-:8])+$signed(-{in[1143-:8],2'b0})+$signed({in[1151-:8],1'b0})+$signed(sharing24)+$signed(-1);
assign weighted_sum[366] = $signed(-{in[1159-:8],2'b0})+$signed({in[1167-:8],1'b0})+$signed({in[1175-:8],1'b0})+$signed(in[1175-:8])+$signed(-{in[1383-:8],3'b0})+$signed(-{in[1391-:8],3'b0})+$signed({in[943-:8],1'b0})+$signed({in[951-:8],2'b0})+$signed(-{in[1399-:8],1'b0})+$signed(in[951-:8])+$signed(sharing25)+$signed(-1);
assign weighted_sum[367] = $signed({in[967-:8],2'b0})+$signed(-{in[1415-:8],1'b0})+$signed(in[967-:8])+$signed(-{in[1175-:8],2'b0})+$signed({in[1183-:8],1'b0})+$signed({in[1191-:8],1'b0})+$signed(in[1191-:8])+$signed(-{in[1399-:8],3'b0})+$signed(-{in[1407-:8],3'b0})+$signed({in[959-:8],1'b0})+$signed(sharing26)+$signed(-1);
assign weighted_sum[368] = $signed(-{in[1415-:8],3'b0})+$signed(-{in[1423-:8],3'b0})+$signed({in[975-:8],1'b0})+$signed({in[983-:8],2'b0})+$signed(-{in[1431-:8],1'b0})+$signed(in[983-:8])+$signed(-{in[1191-:8],2'b0})+$signed({in[1199-:8],1'b0})+$signed({in[1207-:8],1'b0})+$signed(in[1207-:8])+$signed(sharing151)+$signed(-1);
assign weighted_sum[369] = $signed({in[1223-:8],1'b0})+$signed(in[1223-:8])+$signed(-{in[1431-:8],3'b0})+$signed(-{in[1439-:8],3'b0})+$signed({in[991-:8],1'b0})+$signed({in[999-:8],2'b0})+$signed(-{in[1447-:8],1'b0})+$signed(in[999-:8])+$signed(-{in[1207-:8],2'b0})+$signed({in[1215-:8],1'b0})+$signed(sharing27)+$signed(-1);
assign weighted_sum[370] = $signed(-{in[1223-:8],2'b0})+$signed({in[1231-:8],1'b0})+$signed({in[1239-:8],1'b0})+$signed(in[1239-:8])+$signed(-{in[1447-:8],3'b0})+$signed(-{in[1455-:8],3'b0})+$signed({in[1007-:8],1'b0})+$signed({in[1015-:8],2'b0})+$signed(-{in[1463-:8],1'b0})+$signed(in[1015-:8])+$signed(sharing28)+$signed(-1);
assign weighted_sum[371] = $signed({in[1031-:8],2'b0})+$signed(-{in[1479-:8],1'b0})+$signed(in[1031-:8])+$signed(-{in[1239-:8],2'b0})+$signed({in[1247-:8],1'b0})+$signed({in[1255-:8],1'b0})+$signed(in[1255-:8])+$signed(-{in[1463-:8],3'b0})+$signed(-{in[1471-:8],3'b0})+$signed({in[1023-:8],1'b0})+$signed(sharing29)+$signed(-1);
assign weighted_sum[372] = $signed(-{in[1479-:8],3'b0})+$signed(-{in[1487-:8],3'b0})+$signed({in[1039-:8],1'b0})+$signed({in[1047-:8],2'b0})+$signed(-{in[1495-:8],1'b0})+$signed(in[1047-:8])+$signed(-{in[1255-:8],2'b0})+$signed({in[1263-:8],1'b0})+$signed({in[1271-:8],1'b0})+$signed(in[1271-:8])+$signed(sharing30)+$signed(-1);
assign weighted_sum[373] = $signed({in[1287-:8],1'b0})+$signed(in[1287-:8])+$signed(-{in[1495-:8],3'b0})+$signed(-{in[1503-:8],3'b0})+$signed({in[1055-:8],1'b0})+$signed({in[1063-:8],2'b0})+$signed(-{in[1511-:8],1'b0})+$signed(in[1063-:8])+$signed(-{in[1271-:8],2'b0})+$signed({in[1279-:8],1'b0})+$signed(sharing31)+$signed(-1);
assign weighted_sum[374] = $signed(-{in[1287-:8],2'b0})+$signed({in[1295-:8],1'b0})+$signed({in[1303-:8],1'b0})+$signed(in[1303-:8])+$signed(-{in[1511-:8],3'b0})+$signed(-{in[1519-:8],3'b0})+$signed({in[1071-:8],1'b0})+$signed({in[1079-:8],2'b0})+$signed(-{in[1527-:8],1'b0})+$signed(in[1079-:8])+$signed(sharing32)+$signed(-1);
assign weighted_sum[375] = $signed({in[1095-:8],2'b0})+$signed(-{in[1543-:8],1'b0})+$signed(in[1095-:8])+$signed(-{in[1303-:8],2'b0})+$signed({in[1311-:8],1'b0})+$signed({in[1319-:8],1'b0})+$signed(in[1319-:8])+$signed(-{in[1527-:8],3'b0})+$signed(-{in[1535-:8],3'b0})+$signed({in[1087-:8],1'b0})+$signed(sharing33)+$signed(-1);
assign weighted_sum[376] = $signed(-{in[1543-:8],3'b0})+$signed(-{in[1551-:8],3'b0})+$signed({in[1103-:8],1'b0})+$signed({in[1111-:8],2'b0})+$signed(-{in[1559-:8],1'b0})+$signed(in[1111-:8])+$signed(-{in[1319-:8],2'b0})+$signed({in[1327-:8],1'b0})+$signed({in[1335-:8],1'b0})+$signed(in[1335-:8])+$signed(sharing152)+$signed(-1);
assign weighted_sum[377] = $signed(-{in[1799-:8],3'b0})+$signed(-{in[1807-:8],3'b0})+$signed({in[1359-:8],1'b0})+$signed({in[1367-:8],2'b0})+$signed(-{in[1815-:8],1'b0})+$signed(in[1367-:8])+$signed(-{in[1575-:8],2'b0})+$signed({in[1583-:8],1'b0})+$signed({in[1591-:8],1'b0})+$signed(in[1591-:8])+$signed(sharing34)+$signed(-1);
assign weighted_sum[378] = $signed({in[1607-:8],1'b0})+$signed(in[1607-:8])+$signed(-{in[1815-:8],3'b0})+$signed(-{in[1823-:8],3'b0})+$signed({in[1375-:8],1'b0})+$signed({in[1383-:8],2'b0})+$signed(-{in[1831-:8],1'b0})+$signed(in[1383-:8])+$signed(-{in[1591-:8],2'b0})+$signed({in[1599-:8],1'b0})+$signed(sharing35)+$signed(-1);
assign weighted_sum[379] = $signed(-{in[1607-:8],2'b0})+$signed({in[1615-:8],1'b0})+$signed({in[1623-:8],1'b0})+$signed(in[1623-:8])+$signed(-{in[1831-:8],3'b0})+$signed(-{in[1839-:8],3'b0})+$signed({in[1391-:8],1'b0})+$signed({in[1399-:8],2'b0})+$signed(-{in[1847-:8],1'b0})+$signed(in[1399-:8])+$signed(sharing36)+$signed(-1);
assign weighted_sum[380] = $signed({in[1415-:8],2'b0})+$signed(-{in[1863-:8],1'b0})+$signed(in[1415-:8])+$signed(-{in[1623-:8],2'b0})+$signed({in[1631-:8],1'b0})+$signed({in[1639-:8],1'b0})+$signed(in[1639-:8])+$signed(-{in[1847-:8],3'b0})+$signed(-{in[1855-:8],3'b0})+$signed({in[1407-:8],1'b0})+$signed(sharing37)+$signed(-1);
assign weighted_sum[381] = $signed(-{in[1863-:8],3'b0})+$signed(-{in[1871-:8],3'b0})+$signed({in[1423-:8],1'b0})+$signed({in[1431-:8],2'b0})+$signed(-{in[1879-:8],1'b0})+$signed(in[1431-:8])+$signed(-{in[1639-:8],2'b0})+$signed({in[1647-:8],1'b0})+$signed({in[1655-:8],1'b0})+$signed(in[1655-:8])+$signed(sharing38)+$signed(-1);
assign weighted_sum[382] = $signed({in[1671-:8],1'b0})+$signed(in[1671-:8])+$signed(-{in[1879-:8],3'b0})+$signed(-{in[1887-:8],3'b0})+$signed({in[1439-:8],1'b0})+$signed({in[1447-:8],2'b0})+$signed(-{in[1895-:8],1'b0})+$signed(in[1447-:8])+$signed(-{in[1655-:8],2'b0})+$signed({in[1663-:8],1'b0})+$signed(sharing39)+$signed(-1);
assign weighted_sum[383] = $signed(-{in[1671-:8],2'b0})+$signed({in[1679-:8],1'b0})+$signed({in[1687-:8],1'b0})+$signed(in[1687-:8])+$signed(-{in[1895-:8],3'b0})+$signed(-{in[1903-:8],3'b0})+$signed({in[1455-:8],1'b0})+$signed({in[1463-:8],2'b0})+$signed(-{in[1911-:8],1'b0})+$signed(in[1463-:8])+$signed(sharing40)+$signed(-1);
assign weighted_sum[384] = $signed({in[1479-:8],2'b0})+$signed(-{in[1927-:8],1'b0})+$signed(in[1479-:8])+$signed(-{in[1687-:8],2'b0})+$signed({in[1695-:8],1'b0})+$signed({in[1703-:8],1'b0})+$signed(in[1703-:8])+$signed(-{in[1911-:8],3'b0})+$signed(-{in[1919-:8],3'b0})+$signed({in[1471-:8],1'b0})+$signed(sharing153)+$signed(-1);
assign weighted_sum[385] = $signed(-{in[1927-:8],3'b0})+$signed(-{in[1935-:8],3'b0})+$signed({in[1487-:8],1'b0})+$signed({in[1495-:8],2'b0})+$signed(-{in[1943-:8],1'b0})+$signed(in[1495-:8])+$signed(-{in[1703-:8],2'b0})+$signed({in[1711-:8],1'b0})+$signed({in[1719-:8],1'b0})+$signed(in[1719-:8])+$signed(sharing41)+$signed(-1);
assign weighted_sum[386] = $signed({in[1735-:8],1'b0})+$signed(in[1735-:8])+$signed(-{in[1943-:8],3'b0})+$signed(-{in[1951-:8],3'b0})+$signed({in[1503-:8],1'b0})+$signed({in[1511-:8],2'b0})+$signed(-{in[1959-:8],1'b0})+$signed(in[1511-:8])+$signed(-{in[1719-:8],2'b0})+$signed({in[1727-:8],1'b0})+$signed(sharing42)+$signed(-1);
assign weighted_sum[387] = $signed(-{in[1735-:8],2'b0})+$signed({in[1743-:8],1'b0})+$signed({in[1751-:8],1'b0})+$signed(in[1751-:8])+$signed(-{in[1959-:8],3'b0})+$signed(-{in[1967-:8],3'b0})+$signed({in[1519-:8],1'b0})+$signed({in[1527-:8],2'b0})+$signed(-{in[1975-:8],1'b0})+$signed(in[1527-:8])+$signed(sharing43)+$signed(-1);
assign weighted_sum[388] = $signed({in[1543-:8],2'b0})+$signed(-{in[1991-:8],1'b0})+$signed(in[1543-:8])+$signed(-{in[1751-:8],2'b0})+$signed({in[1759-:8],1'b0})+$signed({in[1767-:8],1'b0})+$signed(in[1767-:8])+$signed(-{in[1975-:8],3'b0})+$signed(-{in[1983-:8],3'b0})+$signed({in[1535-:8],1'b0})+$signed(sharing44)+$signed(-1);
assign weighted_sum[389] = $signed(-{in[1991-:8],3'b0})+$signed(-{in[1999-:8],3'b0})+$signed({in[1551-:8],1'b0})+$signed({in[1559-:8],2'b0})+$signed(-{in[2007-:8],1'b0})+$signed(in[1559-:8])+$signed(-{in[1767-:8],2'b0})+$signed({in[1775-:8],1'b0})+$signed({in[1783-:8],1'b0})+$signed(in[1783-:8])+$signed(sharing45)+$signed(-1);
assign weighted_sum[390] = $signed(-{in[2247-:8],3'b0})+$signed(-{in[2255-:8],3'b0})+$signed({in[1807-:8],1'b0})+$signed({in[1815-:8],2'b0})+$signed(-{in[2263-:8],1'b0})+$signed(in[1815-:8])+$signed(-{in[2023-:8],2'b0})+$signed({in[2031-:8],1'b0})+$signed({in[2039-:8],1'b0})+$signed(in[2039-:8])+$signed(sharing46)+$signed(-1);
assign weighted_sum[391] = $signed({in[2055-:8],1'b0})+$signed(in[2055-:8])+$signed(-{in[2263-:8],3'b0})+$signed(-{in[2271-:8],3'b0})+$signed({in[1823-:8],1'b0})+$signed({in[1831-:8],2'b0})+$signed(-{in[2279-:8],1'b0})+$signed(in[1831-:8])+$signed(-{in[2039-:8],2'b0})+$signed({in[2047-:8],1'b0})+$signed(sharing47)+$signed(-1);
assign weighted_sum[392] = $signed(-{in[2055-:8],2'b0})+$signed({in[2063-:8],1'b0})+$signed({in[2071-:8],1'b0})+$signed(in[2071-:8])+$signed(-{in[2279-:8],3'b0})+$signed(-{in[2287-:8],3'b0})+$signed({in[1839-:8],1'b0})+$signed({in[1847-:8],2'b0})+$signed(-{in[2295-:8],1'b0})+$signed(in[1847-:8])+$signed(sharing154)+$signed(-1);
assign weighted_sum[393] = $signed({in[1863-:8],2'b0})+$signed(-{in[2311-:8],1'b0})+$signed(in[1863-:8])+$signed(-{in[2071-:8],2'b0})+$signed({in[2079-:8],1'b0})+$signed({in[2087-:8],1'b0})+$signed(in[2087-:8])+$signed(-{in[2295-:8],3'b0})+$signed(-{in[2303-:8],3'b0})+$signed({in[1855-:8],1'b0})+$signed(sharing48)+$signed(-1);
assign weighted_sum[394] = $signed(-{in[2311-:8],3'b0})+$signed(-{in[2319-:8],3'b0})+$signed({in[1871-:8],1'b0})+$signed({in[1879-:8],2'b0})+$signed(-{in[2327-:8],1'b0})+$signed(in[1879-:8])+$signed(-{in[2087-:8],2'b0})+$signed({in[2095-:8],1'b0})+$signed({in[2103-:8],1'b0})+$signed(in[2103-:8])+$signed(sharing49)+$signed(-1);
assign weighted_sum[395] = $signed({in[2119-:8],1'b0})+$signed(in[2119-:8])+$signed(-{in[2327-:8],3'b0})+$signed(-{in[2335-:8],3'b0})+$signed({in[1887-:8],1'b0})+$signed({in[1895-:8],2'b0})+$signed(-{in[2343-:8],1'b0})+$signed(in[1895-:8])+$signed(-{in[2103-:8],2'b0})+$signed({in[2111-:8],1'b0})+$signed(sharing50)+$signed(-1);
assign weighted_sum[396] = $signed(-{in[2119-:8],2'b0})+$signed({in[2127-:8],1'b0})+$signed({in[2135-:8],1'b0})+$signed(in[2135-:8])+$signed(-{in[2343-:8],3'b0})+$signed(-{in[2351-:8],3'b0})+$signed({in[1903-:8],1'b0})+$signed({in[1911-:8],2'b0})+$signed(-{in[2359-:8],1'b0})+$signed(in[1911-:8])+$signed(sharing51)+$signed(-1);
assign weighted_sum[397] = $signed({in[1927-:8],2'b0})+$signed(-{in[2375-:8],1'b0})+$signed(in[1927-:8])+$signed(-{in[2135-:8],2'b0})+$signed({in[2143-:8],1'b0})+$signed({in[2151-:8],1'b0})+$signed(in[2151-:8])+$signed(-{in[2359-:8],3'b0})+$signed(-{in[2367-:8],3'b0})+$signed({in[1919-:8],1'b0})+$signed(sharing52)+$signed(-1);
assign weighted_sum[398] = $signed(-{in[2375-:8],3'b0})+$signed(-{in[2383-:8],3'b0})+$signed({in[1935-:8],1'b0})+$signed({in[1943-:8],2'b0})+$signed(-{in[2391-:8],1'b0})+$signed(in[1943-:8])+$signed(-{in[2151-:8],2'b0})+$signed({in[2159-:8],1'b0})+$signed({in[2167-:8],1'b0})+$signed(in[2167-:8])+$signed(sharing53)+$signed(-1);
assign weighted_sum[399] = $signed({in[2183-:8],1'b0})+$signed(in[2183-:8])+$signed(-{in[2391-:8],3'b0})+$signed(-{in[2399-:8],3'b0})+$signed({in[1951-:8],1'b0})+$signed({in[1959-:8],2'b0})+$signed(-{in[2407-:8],1'b0})+$signed(in[1959-:8])+$signed(-{in[2167-:8],2'b0})+$signed({in[2175-:8],1'b0})+$signed(sharing54)+$signed(-1);
assign weighted_sum[400] = $signed(-{in[2183-:8],2'b0})+$signed({in[2191-:8],1'b0})+$signed({in[2199-:8],1'b0})+$signed(in[2199-:8])+$signed(-{in[2407-:8],3'b0})+$signed(-{in[2415-:8],3'b0})+$signed({in[1967-:8],1'b0})+$signed({in[1975-:8],2'b0})+$signed(-{in[2423-:8],1'b0})+$signed(in[1975-:8])+$signed(sharing155)+$signed(-1);
assign weighted_sum[401] = $signed({in[1991-:8],2'b0})+$signed(-{in[2439-:8],1'b0})+$signed(in[1991-:8])+$signed(-{in[2199-:8],2'b0})+$signed({in[2207-:8],1'b0})+$signed({in[2215-:8],1'b0})+$signed(in[2215-:8])+$signed(-{in[2423-:8],3'b0})+$signed(-{in[2431-:8],3'b0})+$signed({in[1983-:8],1'b0})+$signed(sharing55)+$signed(-1);
assign weighted_sum[402] = $signed(-{in[2439-:8],3'b0})+$signed(-{in[2447-:8],3'b0})+$signed({in[1999-:8],1'b0})+$signed({in[2007-:8],2'b0})+$signed(-{in[2455-:8],1'b0})+$signed(in[2007-:8])+$signed(-{in[2215-:8],2'b0})+$signed({in[2223-:8],1'b0})+$signed({in[2231-:8],1'b0})+$signed(in[2231-:8])+$signed(sharing56)+$signed(-1);
assign weighted_sum[403] = $signed(-{in[2695-:8],3'b0})+$signed(-{in[2703-:8],3'b0})+$signed({in[2255-:8],1'b0})+$signed({in[2263-:8],2'b0})+$signed(-{in[2711-:8],1'b0})+$signed(in[2263-:8])+$signed(-{in[2471-:8],2'b0})+$signed({in[2479-:8],1'b0})+$signed({in[2487-:8],1'b0})+$signed(in[2487-:8])+$signed(sharing57)+$signed(-1);
assign weighted_sum[404] = $signed({in[2503-:8],1'b0})+$signed(in[2503-:8])+$signed(-{in[2711-:8],3'b0})+$signed(-{in[2719-:8],3'b0})+$signed({in[2271-:8],1'b0})+$signed({in[2279-:8],2'b0})+$signed(-{in[2727-:8],1'b0})+$signed(in[2279-:8])+$signed(-{in[2487-:8],2'b0})+$signed({in[2495-:8],1'b0})+$signed(sharing58)+$signed(-1);
assign weighted_sum[405] = $signed(-{in[2503-:8],2'b0})+$signed({in[2511-:8],1'b0})+$signed({in[2519-:8],1'b0})+$signed(in[2519-:8])+$signed(-{in[2727-:8],3'b0})+$signed(-{in[2735-:8],3'b0})+$signed({in[2287-:8],1'b0})+$signed({in[2295-:8],2'b0})+$signed(-{in[2743-:8],1'b0})+$signed(in[2295-:8])+$signed(sharing59)+$signed(-1);
assign weighted_sum[406] = $signed({in[2311-:8],2'b0})+$signed(-{in[2759-:8],1'b0})+$signed(in[2311-:8])+$signed(-{in[2519-:8],2'b0})+$signed({in[2527-:8],1'b0})+$signed({in[2535-:8],1'b0})+$signed(in[2535-:8])+$signed(-{in[2743-:8],3'b0})+$signed(-{in[2751-:8],3'b0})+$signed({in[2303-:8],1'b0})+$signed(sharing60)+$signed(-1);
assign weighted_sum[407] = $signed(-{in[2759-:8],3'b0})+$signed(-{in[2767-:8],3'b0})+$signed({in[2319-:8],1'b0})+$signed({in[2327-:8],2'b0})+$signed(-{in[2775-:8],1'b0})+$signed(in[2327-:8])+$signed(-{in[2535-:8],2'b0})+$signed({in[2543-:8],1'b0})+$signed({in[2551-:8],1'b0})+$signed(in[2551-:8])+$signed(sharing61)+$signed(-1);
assign weighted_sum[408] = $signed({in[2567-:8],1'b0})+$signed(in[2567-:8])+$signed(-{in[2775-:8],3'b0})+$signed(-{in[2783-:8],3'b0})+$signed({in[2335-:8],1'b0})+$signed({in[2343-:8],2'b0})+$signed(-{in[2791-:8],1'b0})+$signed(in[2343-:8])+$signed(-{in[2551-:8],2'b0})+$signed({in[2559-:8],1'b0})+$signed(sharing156)+$signed(-1);
assign weighted_sum[409] = $signed(-{in[2567-:8],2'b0})+$signed({in[2575-:8],1'b0})+$signed({in[2583-:8],1'b0})+$signed(in[2583-:8])+$signed(-{in[2791-:8],3'b0})+$signed(-{in[2799-:8],3'b0})+$signed({in[2351-:8],1'b0})+$signed({in[2359-:8],2'b0})+$signed(-{in[2807-:8],1'b0})+$signed(in[2359-:8])+$signed(sharing62)+$signed(-1);
assign weighted_sum[410] = $signed({in[2375-:8],2'b0})+$signed(-{in[2823-:8],1'b0})+$signed(in[2375-:8])+$signed(-{in[2583-:8],2'b0})+$signed({in[2591-:8],1'b0})+$signed({in[2599-:8],1'b0})+$signed(in[2599-:8])+$signed(-{in[2807-:8],3'b0})+$signed(-{in[2815-:8],3'b0})+$signed({in[2367-:8],1'b0})+$signed(sharing63)+$signed(-1);
assign weighted_sum[411] = $signed(-{in[2823-:8],3'b0})+$signed(-{in[2831-:8],3'b0})+$signed({in[2383-:8],1'b0})+$signed({in[2391-:8],2'b0})+$signed(-{in[2839-:8],1'b0})+$signed(in[2391-:8])+$signed(-{in[2599-:8],2'b0})+$signed({in[2607-:8],1'b0})+$signed({in[2615-:8],1'b0})+$signed(in[2615-:8])+$signed(sharing64)+$signed(-1);
assign weighted_sum[412] = $signed({in[2631-:8],1'b0})+$signed(in[2631-:8])+$signed(-{in[2839-:8],3'b0})+$signed(-{in[2847-:8],3'b0})+$signed({in[2399-:8],1'b0})+$signed({in[2407-:8],2'b0})+$signed(-{in[2855-:8],1'b0})+$signed(in[2407-:8])+$signed(-{in[2615-:8],2'b0})+$signed({in[2623-:8],1'b0})+$signed(sharing65)+$signed(-1);
assign weighted_sum[413] = $signed(-{in[2631-:8],2'b0})+$signed({in[2639-:8],1'b0})+$signed({in[2647-:8],1'b0})+$signed(in[2647-:8])+$signed(-{in[2855-:8],3'b0})+$signed(-{in[2863-:8],3'b0})+$signed({in[2415-:8],1'b0})+$signed({in[2423-:8],2'b0})+$signed(-{in[2871-:8],1'b0})+$signed(in[2423-:8])+$signed(sharing66)+$signed(-1);
assign weighted_sum[414] = $signed({in[2439-:8],2'b0})+$signed(-{in[2887-:8],1'b0})+$signed(in[2439-:8])+$signed(-{in[2647-:8],2'b0})+$signed({in[2655-:8],1'b0})+$signed({in[2663-:8],1'b0})+$signed(in[2663-:8])+$signed(-{in[2871-:8],3'b0})+$signed(-{in[2879-:8],3'b0})+$signed({in[2431-:8],1'b0})+$signed(sharing67)+$signed(-1);
assign weighted_sum[415] = $signed(-{in[2887-:8],3'b0})+$signed(-{in[2895-:8],3'b0})+$signed({in[2447-:8],1'b0})+$signed({in[2455-:8],2'b0})+$signed(-{in[2903-:8],1'b0})+$signed(in[2455-:8])+$signed(-{in[2663-:8],2'b0})+$signed({in[2671-:8],1'b0})+$signed({in[2679-:8],1'b0})+$signed(in[2679-:8])+$signed(sharing68)+$signed(-1);
assign weighted_sum[416] = $signed(-{in[3143-:8],3'b0})+$signed(-{in[3151-:8],3'b0})+$signed({in[2703-:8],1'b0})+$signed({in[2711-:8],2'b0})+$signed(-{in[3159-:8],1'b0})+$signed(in[2711-:8])+$signed(-{in[2919-:8],2'b0})+$signed({in[2927-:8],1'b0})+$signed({in[2935-:8],1'b0})+$signed(in[2935-:8])+$signed(sharing157)+$signed(-1);
assign weighted_sum[417] = $signed({in[2951-:8],1'b0})+$signed(in[2951-:8])+$signed(-{in[3159-:8],3'b0})+$signed(-{in[3167-:8],3'b0})+$signed({in[2719-:8],1'b0})+$signed({in[2727-:8],2'b0})+$signed(-{in[3175-:8],1'b0})+$signed(in[2727-:8])+$signed(-{in[2935-:8],2'b0})+$signed({in[2943-:8],1'b0})+$signed(sharing69)+$signed(-1);
assign weighted_sum[418] = $signed(-{in[2951-:8],2'b0})+$signed({in[2959-:8],1'b0})+$signed({in[2967-:8],1'b0})+$signed(in[2967-:8])+$signed(-{in[3175-:8],3'b0})+$signed(-{in[3183-:8],3'b0})+$signed({in[2735-:8],1'b0})+$signed({in[2743-:8],2'b0})+$signed(-{in[3191-:8],1'b0})+$signed(in[2743-:8])+$signed(sharing70)+$signed(-1);
assign weighted_sum[419] = $signed({in[2759-:8],2'b0})+$signed(-{in[3207-:8],1'b0})+$signed(in[2759-:8])+$signed(-{in[2967-:8],2'b0})+$signed({in[2975-:8],1'b0})+$signed({in[2983-:8],1'b0})+$signed(in[2983-:8])+$signed(-{in[3191-:8],3'b0})+$signed(-{in[3199-:8],3'b0})+$signed({in[2751-:8],1'b0})+$signed(sharing71)+$signed(-1);
assign weighted_sum[420] = $signed(-{in[3207-:8],3'b0})+$signed(-{in[3215-:8],3'b0})+$signed({in[2767-:8],1'b0})+$signed({in[2775-:8],2'b0})+$signed(-{in[3223-:8],1'b0})+$signed(in[2775-:8])+$signed(-{in[2983-:8],2'b0})+$signed({in[2991-:8],1'b0})+$signed({in[2999-:8],1'b0})+$signed(in[2999-:8])+$signed(sharing72)+$signed(-1);
assign weighted_sum[421] = $signed({in[3015-:8],1'b0})+$signed(in[3015-:8])+$signed(-{in[3223-:8],3'b0})+$signed(-{in[3231-:8],3'b0})+$signed({in[2783-:8],1'b0})+$signed({in[2791-:8],2'b0})+$signed(-{in[3239-:8],1'b0})+$signed(in[2791-:8])+$signed(-{in[2999-:8],2'b0})+$signed({in[3007-:8],1'b0})+$signed(sharing73)+$signed(-1);
assign weighted_sum[422] = $signed(-{in[3015-:8],2'b0})+$signed({in[3023-:8],1'b0})+$signed({in[3031-:8],1'b0})+$signed(in[3031-:8])+$signed(-{in[3239-:8],3'b0})+$signed(-{in[3247-:8],3'b0})+$signed({in[2799-:8],1'b0})+$signed({in[2807-:8],2'b0})+$signed(-{in[3255-:8],1'b0})+$signed(in[2807-:8])+$signed(sharing74)+$signed(-1);
assign weighted_sum[423] = $signed({in[2823-:8],2'b0})+$signed(-{in[3271-:8],1'b0})+$signed(in[2823-:8])+$signed(-{in[3031-:8],2'b0})+$signed({in[3039-:8],1'b0})+$signed({in[3047-:8],1'b0})+$signed(in[3047-:8])+$signed(-{in[3255-:8],3'b0})+$signed(-{in[3263-:8],3'b0})+$signed({in[2815-:8],1'b0})+$signed(sharing75)+$signed(-1);
assign weighted_sum[424] = $signed(-{in[3271-:8],3'b0})+$signed(-{in[3279-:8],3'b0})+$signed({in[2831-:8],1'b0})+$signed({in[2839-:8],2'b0})+$signed(-{in[3287-:8],1'b0})+$signed(in[2839-:8])+$signed(-{in[3047-:8],2'b0})+$signed({in[3055-:8],1'b0})+$signed({in[3063-:8],1'b0})+$signed(in[3063-:8])+$signed(sharing158)+$signed(-1);
assign weighted_sum[425] = $signed({in[3079-:8],1'b0})+$signed(in[3079-:8])+$signed(-{in[3287-:8],3'b0})+$signed(-{in[3295-:8],3'b0})+$signed({in[2847-:8],1'b0})+$signed({in[2855-:8],2'b0})+$signed(-{in[3303-:8],1'b0})+$signed(in[2855-:8])+$signed(-{in[3063-:8],2'b0})+$signed({in[3071-:8],1'b0})+$signed(sharing76)+$signed(-1);
assign weighted_sum[426] = $signed(-{in[3079-:8],2'b0})+$signed({in[3087-:8],1'b0})+$signed({in[3095-:8],1'b0})+$signed(in[3095-:8])+$signed(-{in[3303-:8],3'b0})+$signed(-{in[3311-:8],3'b0})+$signed({in[2863-:8],1'b0})+$signed({in[2871-:8],2'b0})+$signed(-{in[3319-:8],1'b0})+$signed(in[2871-:8])+$signed(sharing77)+$signed(-1);
assign weighted_sum[427] = $signed({in[2887-:8],2'b0})+$signed(-{in[3335-:8],1'b0})+$signed(in[2887-:8])+$signed(-{in[3095-:8],2'b0})+$signed({in[3103-:8],1'b0})+$signed({in[3111-:8],1'b0})+$signed(in[3111-:8])+$signed(-{in[3319-:8],3'b0})+$signed(-{in[3327-:8],3'b0})+$signed({in[2879-:8],1'b0})+$signed(sharing78)+$signed(-1);
assign weighted_sum[428] = $signed(-{in[3335-:8],3'b0})+$signed(-{in[3343-:8],3'b0})+$signed({in[2895-:8],1'b0})+$signed({in[2903-:8],2'b0})+$signed(-{in[3351-:8],1'b0})+$signed(in[2903-:8])+$signed(-{in[3111-:8],2'b0})+$signed({in[3119-:8],1'b0})+$signed({in[3127-:8],1'b0})+$signed(in[3127-:8])+$signed(sharing79)+$signed(-1);
assign weighted_sum[429] = $signed(-{in[3591-:8],3'b0})+$signed(-{in[3599-:8],3'b0})+$signed({in[3151-:8],1'b0})+$signed({in[3159-:8],2'b0})+$signed(-{in[3607-:8],1'b0})+$signed(in[3159-:8])+$signed(-{in[3367-:8],2'b0})+$signed({in[3375-:8],1'b0})+$signed({in[3383-:8],1'b0})+$signed(in[3383-:8])+$signed(sharing80)+$signed(-1);
assign weighted_sum[430] = $signed({in[3399-:8],1'b0})+$signed(in[3399-:8])+$signed(-{in[3607-:8],3'b0})+$signed(-{in[3615-:8],3'b0})+$signed({in[3167-:8],1'b0})+$signed({in[3175-:8],2'b0})+$signed(-{in[3623-:8],1'b0})+$signed(in[3175-:8])+$signed(-{in[3383-:8],2'b0})+$signed({in[3391-:8],1'b0})+$signed(sharing81)+$signed(-1);
assign weighted_sum[431] = $signed(-{in[3399-:8],2'b0})+$signed({in[3407-:8],1'b0})+$signed({in[3415-:8],1'b0})+$signed(in[3415-:8])+$signed(-{in[3623-:8],3'b0})+$signed(-{in[3631-:8],3'b0})+$signed({in[3183-:8],1'b0})+$signed({in[3191-:8],2'b0})+$signed(-{in[3639-:8],1'b0})+$signed(in[3191-:8])+$signed(sharing82)+$signed(-1);
assign weighted_sum[432] = $signed({in[3207-:8],2'b0})+$signed(-{in[3655-:8],1'b0})+$signed(in[3207-:8])+$signed(-{in[3415-:8],2'b0})+$signed({in[3423-:8],1'b0})+$signed({in[3431-:8],1'b0})+$signed(in[3431-:8])+$signed(-{in[3639-:8],3'b0})+$signed(-{in[3647-:8],3'b0})+$signed({in[3199-:8],1'b0})+$signed(sharing159)+$signed(-1);
assign weighted_sum[433] = $signed(-{in[3655-:8],3'b0})+$signed(-{in[3663-:8],3'b0})+$signed({in[3215-:8],1'b0})+$signed({in[3223-:8],2'b0})+$signed(-{in[3671-:8],1'b0})+$signed(in[3223-:8])+$signed(-{in[3431-:8],2'b0})+$signed({in[3439-:8],1'b0})+$signed({in[3447-:8],1'b0})+$signed(in[3447-:8])+$signed(sharing83)+$signed(-1);
assign weighted_sum[434] = $signed({in[3463-:8],1'b0})+$signed(in[3463-:8])+$signed(-{in[3671-:8],3'b0})+$signed(-{in[3679-:8],3'b0})+$signed({in[3231-:8],1'b0})+$signed({in[3239-:8],2'b0})+$signed(-{in[3687-:8],1'b0})+$signed(in[3239-:8])+$signed(-{in[3447-:8],2'b0})+$signed({in[3455-:8],1'b0})+$signed(sharing84)+$signed(-1);
assign weighted_sum[435] = $signed(-{in[3463-:8],2'b0})+$signed({in[3471-:8],1'b0})+$signed({in[3479-:8],1'b0})+$signed(in[3479-:8])+$signed(-{in[3687-:8],3'b0})+$signed(-{in[3695-:8],3'b0})+$signed({in[3247-:8],1'b0})+$signed({in[3255-:8],2'b0})+$signed(-{in[3703-:8],1'b0})+$signed(in[3255-:8])+$signed(sharing85)+$signed(-1);
assign weighted_sum[436] = $signed({in[3271-:8],2'b0})+$signed(-{in[3719-:8],1'b0})+$signed(in[3271-:8])+$signed(-{in[3479-:8],2'b0})+$signed({in[3487-:8],1'b0})+$signed({in[3495-:8],1'b0})+$signed(in[3495-:8])+$signed(-{in[3703-:8],3'b0})+$signed(-{in[3711-:8],3'b0})+$signed({in[3263-:8],1'b0})+$signed(sharing86)+$signed(-1);
assign weighted_sum[437] = $signed(-{in[3719-:8],3'b0})+$signed(-{in[3727-:8],3'b0})+$signed({in[3279-:8],1'b0})+$signed({in[3287-:8],2'b0})+$signed(-{in[3735-:8],1'b0})+$signed(in[3287-:8])+$signed(-{in[3495-:8],2'b0})+$signed({in[3503-:8],1'b0})+$signed({in[3511-:8],1'b0})+$signed(in[3511-:8])+$signed(sharing87)+$signed(-1);
assign weighted_sum[438] = $signed({in[3527-:8],1'b0})+$signed(in[3527-:8])+$signed(-{in[3735-:8],3'b0})+$signed(-{in[3743-:8],3'b0})+$signed({in[3295-:8],1'b0})+$signed({in[3303-:8],2'b0})+$signed(-{in[3751-:8],1'b0})+$signed(in[3303-:8])+$signed(-{in[3511-:8],2'b0})+$signed({in[3519-:8],1'b0})+$signed(sharing88)+$signed(-1);
assign weighted_sum[439] = $signed(-{in[3527-:8],2'b0})+$signed({in[3535-:8],1'b0})+$signed({in[3543-:8],1'b0})+$signed(in[3543-:8])+$signed(-{in[3751-:8],3'b0})+$signed(-{in[3759-:8],3'b0})+$signed({in[3311-:8],1'b0})+$signed({in[3319-:8],2'b0})+$signed(-{in[3767-:8],1'b0})+$signed(in[3319-:8])+$signed(sharing89)+$signed(-1);
assign weighted_sum[440] = $signed({in[3335-:8],2'b0})+$signed(-{in[3783-:8],1'b0})+$signed(in[3335-:8])+$signed(-{in[3543-:8],2'b0})+$signed({in[3551-:8],1'b0})+$signed({in[3559-:8],1'b0})+$signed(in[3559-:8])+$signed(-{in[3767-:8],3'b0})+$signed(-{in[3775-:8],3'b0})+$signed({in[3327-:8],1'b0})+$signed(sharing160)+$signed(-1);
assign weighted_sum[441] = $signed(-{in[3783-:8],3'b0})+$signed(-{in[3791-:8],3'b0})+$signed({in[3343-:8],1'b0})+$signed({in[3351-:8],2'b0})+$signed(-{in[3799-:8],1'b0})+$signed(in[3351-:8])+$signed(-{in[3559-:8],2'b0})+$signed({in[3567-:8],1'b0})+$signed({in[3575-:8],1'b0})+$signed(in[3575-:8])+$signed(sharing90)+$signed(-1);
assign weighted_sum[442] = $signed(-{in[4039-:8],3'b0})+$signed(-{in[4047-:8],3'b0})+$signed({in[3599-:8],1'b0})+$signed({in[3607-:8],2'b0})+$signed(-{in[4055-:8],1'b0})+$signed(in[3607-:8])+$signed(-{in[3815-:8],2'b0})+$signed({in[3823-:8],1'b0})+$signed({in[3831-:8],1'b0})+$signed(in[3831-:8])+$signed(sharing91)+$signed(-1);
assign weighted_sum[443] = $signed({in[3847-:8],1'b0})+$signed(in[3847-:8])+$signed(-{in[4055-:8],3'b0})+$signed(-{in[4063-:8],3'b0})+$signed({in[3615-:8],1'b0})+$signed({in[3623-:8],2'b0})+$signed(-{in[4071-:8],1'b0})+$signed(in[3623-:8])+$signed(-{in[3831-:8],2'b0})+$signed({in[3839-:8],1'b0})+$signed(sharing92)+$signed(-1);
assign weighted_sum[444] = $signed(-{in[3847-:8],2'b0})+$signed({in[3855-:8],1'b0})+$signed({in[3863-:8],1'b0})+$signed(in[3863-:8])+$signed(-{in[4071-:8],3'b0})+$signed(-{in[4079-:8],3'b0})+$signed({in[3631-:8],1'b0})+$signed({in[3639-:8],2'b0})+$signed(-{in[4087-:8],1'b0})+$signed(in[3639-:8])+$signed(sharing93)+$signed(-1);
assign weighted_sum[445] = $signed({in[3655-:8],2'b0})+$signed(-{in[4103-:8],1'b0})+$signed(in[3655-:8])+$signed(-{in[3863-:8],2'b0})+$signed({in[3871-:8],1'b0})+$signed({in[3879-:8],1'b0})+$signed(in[3879-:8])+$signed(-{in[4087-:8],3'b0})+$signed(-{in[4095-:8],3'b0})+$signed({in[3647-:8],1'b0})+$signed(sharing94)+$signed(-1);
assign weighted_sum[446] = $signed(-{in[4103-:8],3'b0})+$signed(-{in[4111-:8],3'b0})+$signed({in[3663-:8],1'b0})+$signed({in[3671-:8],2'b0})+$signed(-{in[4119-:8],1'b0})+$signed(in[3671-:8])+$signed(-{in[3879-:8],2'b0})+$signed({in[3887-:8],1'b0})+$signed({in[3895-:8],1'b0})+$signed(in[3895-:8])+$signed(sharing95)+$signed(-1);
assign weighted_sum[447] = $signed({in[3911-:8],1'b0})+$signed(in[3911-:8])+$signed(-{in[4119-:8],3'b0})+$signed(-{in[4127-:8],3'b0})+$signed({in[3679-:8],1'b0})+$signed({in[3687-:8],2'b0})+$signed(-{in[4135-:8],1'b0})+$signed(in[3687-:8])+$signed(-{in[3895-:8],2'b0})+$signed({in[3903-:8],1'b0})+$signed(sharing96)+$signed(-1);
assign weighted_sum[448] = $signed(-{in[3911-:8],2'b0})+$signed({in[3919-:8],1'b0})+$signed({in[3927-:8],1'b0})+$signed(in[3927-:8])+$signed(-{in[4135-:8],3'b0})+$signed(-{in[4143-:8],3'b0})+$signed({in[3695-:8],1'b0})+$signed({in[3703-:8],2'b0})+$signed(-{in[4151-:8],1'b0})+$signed(in[3703-:8])+$signed(sharing161)+$signed(-1);
assign weighted_sum[449] = $signed({in[3719-:8],2'b0})+$signed(-{in[4167-:8],1'b0})+$signed(in[3719-:8])+$signed(-{in[3927-:8],2'b0})+$signed({in[3935-:8],1'b0})+$signed({in[3943-:8],1'b0})+$signed(in[3943-:8])+$signed(-{in[4151-:8],3'b0})+$signed(-{in[4159-:8],3'b0})+$signed({in[3711-:8],1'b0})+$signed(sharing97)+$signed(-1);
assign weighted_sum[450] = $signed(-{in[4167-:8],3'b0})+$signed(-{in[4175-:8],3'b0})+$signed({in[3727-:8],1'b0})+$signed({in[3735-:8],2'b0})+$signed(-{in[4183-:8],1'b0})+$signed(in[3735-:8])+$signed(-{in[3943-:8],2'b0})+$signed({in[3951-:8],1'b0})+$signed({in[3959-:8],1'b0})+$signed(in[3959-:8])+$signed(sharing98)+$signed(-1);
assign weighted_sum[451] = $signed({in[3975-:8],1'b0})+$signed(in[3975-:8])+$signed(-{in[4183-:8],3'b0})+$signed(-{in[4191-:8],3'b0})+$signed({in[3743-:8],1'b0})+$signed({in[3751-:8],2'b0})+$signed(-{in[4199-:8],1'b0})+$signed(in[3751-:8])+$signed(-{in[3959-:8],2'b0})+$signed({in[3967-:8],1'b0})+$signed(sharing99)+$signed(-1);
assign weighted_sum[452] = $signed(-{in[3975-:8],2'b0})+$signed({in[3983-:8],1'b0})+$signed({in[3991-:8],1'b0})+$signed(in[3991-:8])+$signed(-{in[4199-:8],3'b0})+$signed(-{in[4207-:8],3'b0})+$signed({in[3759-:8],1'b0})+$signed({in[3767-:8],2'b0})+$signed(-{in[4215-:8],1'b0})+$signed(in[3767-:8])+$signed(sharing100)+$signed(-1);
assign weighted_sum[453] = $signed({in[3783-:8],2'b0})+$signed(-{in[4231-:8],1'b0})+$signed(in[3783-:8])+$signed(-{in[3991-:8],2'b0})+$signed({in[3999-:8],1'b0})+$signed({in[4007-:8],1'b0})+$signed(in[4007-:8])+$signed(-{in[4215-:8],3'b0})+$signed(-{in[4223-:8],3'b0})+$signed({in[3775-:8],1'b0})+$signed(sharing101)+$signed(-1);
assign weighted_sum[454] = $signed(-{in[4231-:8],3'b0})+$signed(-{in[4239-:8],3'b0})+$signed({in[3791-:8],1'b0})+$signed({in[3799-:8],2'b0})+$signed(-{in[4247-:8],1'b0})+$signed(in[3799-:8])+$signed(-{in[4007-:8],2'b0})+$signed({in[4015-:8],1'b0})+$signed({in[4023-:8],1'b0})+$signed(in[4023-:8])+$signed(sharing102)+$signed(-1);
assign weighted_sum[455] = $signed(-{in[4487-:8],3'b0})+$signed(-{in[4495-:8],3'b0})+$signed({in[4047-:8],1'b0})+$signed({in[4055-:8],2'b0})+$signed(-{in[4503-:8],1'b0})+$signed(in[4055-:8])+$signed(-{in[4263-:8],2'b0})+$signed({in[4271-:8],1'b0})+$signed({in[4279-:8],1'b0})+$signed(in[4279-:8])+$signed(sharing103)+$signed(-1);
assign weighted_sum[456] = $signed({in[4295-:8],1'b0})+$signed(in[4295-:8])+$signed(-{in[4503-:8],3'b0})+$signed(-{in[4511-:8],3'b0})+$signed({in[4063-:8],1'b0})+$signed({in[4071-:8],2'b0})+$signed(-{in[4519-:8],1'b0})+$signed(in[4071-:8])+$signed(-{in[4279-:8],2'b0})+$signed({in[4287-:8],1'b0})+$signed(sharing162)+$signed(-1);
assign weighted_sum[457] = $signed(-{in[4295-:8],2'b0})+$signed({in[4303-:8],1'b0})+$signed({in[4311-:8],1'b0})+$signed(in[4311-:8])+$signed(-{in[4519-:8],3'b0})+$signed(-{in[4527-:8],3'b0})+$signed({in[4079-:8],1'b0})+$signed({in[4087-:8],2'b0})+$signed(-{in[4535-:8],1'b0})+$signed(in[4087-:8])+$signed(sharing104)+$signed(-1);
assign weighted_sum[458] = $signed({in[4103-:8],2'b0})+$signed(-{in[4551-:8],1'b0})+$signed(in[4103-:8])+$signed(-{in[4311-:8],2'b0})+$signed({in[4319-:8],1'b0})+$signed({in[4327-:8],1'b0})+$signed(in[4327-:8])+$signed(-{in[4535-:8],3'b0})+$signed(-{in[4543-:8],3'b0})+$signed({in[4095-:8],1'b0})+$signed(sharing105)+$signed(-1);
assign weighted_sum[459] = $signed(-{in[4551-:8],3'b0})+$signed(-{in[4559-:8],3'b0})+$signed({in[4111-:8],1'b0})+$signed({in[4119-:8],2'b0})+$signed(-{in[4567-:8],1'b0})+$signed(in[4119-:8])+$signed(-{in[4327-:8],2'b0})+$signed({in[4335-:8],1'b0})+$signed({in[4343-:8],1'b0})+$signed(in[4343-:8])+$signed(sharing106)+$signed(-1);
assign weighted_sum[460] = $signed({in[4359-:8],1'b0})+$signed(in[4359-:8])+$signed(-{in[4567-:8],3'b0})+$signed(-{in[4575-:8],3'b0})+$signed({in[4127-:8],1'b0})+$signed({in[4135-:8],2'b0})+$signed(-{in[4583-:8],1'b0})+$signed(in[4135-:8])+$signed(-{in[4343-:8],2'b0})+$signed({in[4351-:8],1'b0})+$signed(sharing107)+$signed(-1);
assign weighted_sum[461] = $signed(-{in[4359-:8],2'b0})+$signed({in[4367-:8],1'b0})+$signed({in[4375-:8],1'b0})+$signed(in[4375-:8])+$signed(-{in[4583-:8],3'b0})+$signed(-{in[4591-:8],3'b0})+$signed({in[4143-:8],1'b0})+$signed({in[4151-:8],2'b0})+$signed(-{in[4599-:8],1'b0})+$signed(in[4151-:8])+$signed(sharing108)+$signed(-1);
assign weighted_sum[462] = $signed({in[4167-:8],2'b0})+$signed(-{in[4615-:8],1'b0})+$signed(in[4167-:8])+$signed(-{in[4375-:8],2'b0})+$signed({in[4383-:8],1'b0})+$signed({in[4391-:8],1'b0})+$signed(in[4391-:8])+$signed(-{in[4599-:8],3'b0})+$signed(-{in[4607-:8],3'b0})+$signed({in[4159-:8],1'b0})+$signed(sharing109)+$signed(-1);
assign weighted_sum[463] = $signed(-{in[4615-:8],3'b0})+$signed(-{in[4623-:8],3'b0})+$signed({in[4175-:8],1'b0})+$signed({in[4183-:8],2'b0})+$signed(-{in[4631-:8],1'b0})+$signed(in[4183-:8])+$signed(-{in[4391-:8],2'b0})+$signed({in[4399-:8],1'b0})+$signed({in[4407-:8],1'b0})+$signed(in[4407-:8])+$signed(sharing110)+$signed(-1);
assign weighted_sum[464] = $signed({in[4423-:8],1'b0})+$signed(in[4423-:8])+$signed(-{in[4631-:8],3'b0})+$signed(-{in[4639-:8],3'b0})+$signed({in[4191-:8],1'b0})+$signed({in[4199-:8],2'b0})+$signed(-{in[4647-:8],1'b0})+$signed(in[4199-:8])+$signed(-{in[4407-:8],2'b0})+$signed({in[4415-:8],1'b0})+$signed(sharing163)+$signed(-1);
assign weighted_sum[465] = $signed(-{in[4423-:8],2'b0})+$signed({in[4431-:8],1'b0})+$signed({in[4439-:8],1'b0})+$signed(in[4439-:8])+$signed(-{in[4647-:8],3'b0})+$signed(-{in[4655-:8],3'b0})+$signed({in[4207-:8],1'b0})+$signed({in[4215-:8],2'b0})+$signed(-{in[4663-:8],1'b0})+$signed(in[4215-:8])+$signed(sharing111)+$signed(-1);
assign weighted_sum[466] = $signed({in[4231-:8],2'b0})+$signed(-{in[4679-:8],1'b0})+$signed(in[4231-:8])+$signed(-{in[4439-:8],2'b0})+$signed({in[4447-:8],1'b0})+$signed({in[4455-:8],1'b0})+$signed(in[4455-:8])+$signed(-{in[4663-:8],3'b0})+$signed(-{in[4671-:8],3'b0})+$signed({in[4223-:8],1'b0})+$signed(sharing112)+$signed(-1);
assign weighted_sum[467] = $signed(-{in[4679-:8],3'b0})+$signed(-{in[4687-:8],3'b0})+$signed({in[4239-:8],1'b0})+$signed({in[4247-:8],2'b0})+$signed(-{in[4695-:8],1'b0})+$signed(in[4247-:8])+$signed(-{in[4455-:8],2'b0})+$signed({in[4463-:8],1'b0})+$signed({in[4471-:8],1'b0})+$signed(in[4471-:8])+$signed(sharing113)+$signed(-1);
assign weighted_sum[468] = $signed(-{in[4935-:8],3'b0})+$signed(-{in[4943-:8],3'b0})+$signed({in[4495-:8],1'b0})+$signed({in[4503-:8],2'b0})+$signed(-{in[4951-:8],1'b0})+$signed(in[4503-:8])+$signed(-{in[4711-:8],2'b0})+$signed({in[4719-:8],1'b0})+$signed({in[4727-:8],1'b0})+$signed(in[4727-:8])+$signed(sharing114)+$signed(-1);
assign weighted_sum[469] = $signed({in[4743-:8],1'b0})+$signed(in[4743-:8])+$signed(-{in[4951-:8],3'b0})+$signed(-{in[4959-:8],3'b0})+$signed({in[4511-:8],1'b0})+$signed({in[4519-:8],2'b0})+$signed(-{in[4967-:8],1'b0})+$signed(in[4519-:8])+$signed(-{in[4727-:8],2'b0})+$signed({in[4735-:8],1'b0})+$signed(sharing115)+$signed(-1);
assign weighted_sum[470] = $signed(-{in[4743-:8],2'b0})+$signed({in[4751-:8],1'b0})+$signed({in[4759-:8],1'b0})+$signed(in[4759-:8])+$signed(-{in[4967-:8],3'b0})+$signed(-{in[4975-:8],3'b0})+$signed({in[4527-:8],1'b0})+$signed({in[4535-:8],2'b0})+$signed(-{in[4983-:8],1'b0})+$signed(in[4535-:8])+$signed(sharing116)+$signed(-1);
assign weighted_sum[471] = $signed({in[4551-:8],2'b0})+$signed(-{in[4999-:8],1'b0})+$signed(in[4551-:8])+$signed(-{in[4759-:8],2'b0})+$signed({in[4767-:8],1'b0})+$signed({in[4775-:8],1'b0})+$signed(in[4775-:8])+$signed(-{in[4983-:8],3'b0})+$signed(-{in[4991-:8],3'b0})+$signed({in[4543-:8],1'b0})+$signed(sharing117)+$signed(-1);
assign weighted_sum[472] = $signed(-{in[4999-:8],3'b0})+$signed(-{in[5007-:8],3'b0})+$signed({in[4559-:8],1'b0})+$signed({in[4567-:8],2'b0})+$signed(-{in[5015-:8],1'b0})+$signed(in[4567-:8])+$signed(-{in[4775-:8],2'b0})+$signed({in[4783-:8],1'b0})+$signed({in[4791-:8],1'b0})+$signed(in[4791-:8])+$signed(sharing164)+$signed(-1);
assign weighted_sum[473] = $signed({in[4807-:8],1'b0})+$signed(in[4807-:8])+$signed(-{in[5015-:8],3'b0})+$signed(-{in[5023-:8],3'b0})+$signed({in[4575-:8],1'b0})+$signed({in[4583-:8],2'b0})+$signed(-{in[5031-:8],1'b0})+$signed(in[4583-:8])+$signed(-{in[4791-:8],2'b0})+$signed({in[4799-:8],1'b0})+$signed(sharing118)+$signed(-1);
assign weighted_sum[474] = $signed(-{in[4807-:8],2'b0})+$signed({in[4815-:8],1'b0})+$signed({in[4823-:8],1'b0})+$signed(in[4823-:8])+$signed(-{in[5031-:8],3'b0})+$signed(-{in[5039-:8],3'b0})+$signed({in[4591-:8],1'b0})+$signed({in[4599-:8],2'b0})+$signed(-{in[5047-:8],1'b0})+$signed(in[4599-:8])+$signed(sharing119)+$signed(-1);
assign weighted_sum[475] = $signed({in[4615-:8],2'b0})+$signed(-{in[5063-:8],1'b0})+$signed(in[4615-:8])+$signed(-{in[4823-:8],2'b0})+$signed({in[4831-:8],1'b0})+$signed({in[4839-:8],1'b0})+$signed(in[4839-:8])+$signed(-{in[5047-:8],3'b0})+$signed(-{in[5055-:8],3'b0})+$signed({in[4607-:8],1'b0})+$signed(sharing120)+$signed(-1);
assign weighted_sum[476] = $signed(-{in[5063-:8],3'b0})+$signed(-{in[5071-:8],3'b0})+$signed({in[4623-:8],1'b0})+$signed({in[4631-:8],2'b0})+$signed(-{in[5079-:8],1'b0})+$signed(in[4631-:8])+$signed(-{in[4839-:8],2'b0})+$signed({in[4847-:8],1'b0})+$signed({in[4855-:8],1'b0})+$signed(in[4855-:8])+$signed(sharing121)+$signed(-1);
assign weighted_sum[477] = $signed({in[4871-:8],1'b0})+$signed(in[4871-:8])+$signed(-{in[5079-:8],3'b0})+$signed(-{in[5087-:8],3'b0})+$signed({in[4639-:8],1'b0})+$signed({in[4647-:8],2'b0})+$signed(-{in[5095-:8],1'b0})+$signed(in[4647-:8])+$signed(-{in[4855-:8],2'b0})+$signed({in[4863-:8],1'b0})+$signed(sharing122)+$signed(-1);
assign weighted_sum[478] = $signed(-{in[4871-:8],2'b0})+$signed({in[4879-:8],1'b0})+$signed({in[4887-:8],1'b0})+$signed(in[4887-:8])+$signed(-{in[5095-:8],3'b0})+$signed(-{in[5103-:8],3'b0})+$signed({in[4655-:8],1'b0})+$signed({in[4663-:8],2'b0})+$signed(-{in[5111-:8],1'b0})+$signed(in[4663-:8])+$signed(sharing123)+$signed(-1);
assign weighted_sum[479] = $signed({in[4679-:8],2'b0})+$signed(-{in[5127-:8],1'b0})+$signed(in[4679-:8])+$signed(-{in[4887-:8],2'b0})+$signed({in[4895-:8],1'b0})+$signed({in[4903-:8],1'b0})+$signed(in[4903-:8])+$signed(-{in[5111-:8],3'b0})+$signed(-{in[5119-:8],3'b0})+$signed({in[4671-:8],1'b0})+$signed(sharing124)+$signed(-1);
assign weighted_sum[480] = $signed(-{in[5127-:8],3'b0})+$signed(-{in[5135-:8],3'b0})+$signed({in[4687-:8],1'b0})+$signed({in[4695-:8],2'b0})+$signed(-{in[5143-:8],1'b0})+$signed(in[4695-:8])+$signed(-{in[4903-:8],2'b0})+$signed({in[4911-:8],1'b0})+$signed({in[4919-:8],1'b0})+$signed(in[4919-:8])+$signed(sharing165)+$signed(-1);
assign weighted_sum[481] = $signed(-{in[5383-:8],3'b0})+$signed(-{in[5391-:8],3'b0})+$signed({in[4943-:8],1'b0})+$signed({in[4951-:8],2'b0})+$signed(-{in[5399-:8],1'b0})+$signed(in[4951-:8])+$signed(-{in[5159-:8],2'b0})+$signed({in[5167-:8],1'b0})+$signed({in[5175-:8],1'b0})+$signed(in[5175-:8])+$signed(sharing125)+$signed(-1);
assign weighted_sum[482] = $signed({in[5191-:8],1'b0})+$signed(in[5191-:8])+$signed(-{in[5399-:8],3'b0})+$signed(-{in[5407-:8],3'b0})+$signed({in[4959-:8],1'b0})+$signed({in[4967-:8],2'b0})+$signed(-{in[5415-:8],1'b0})+$signed(in[4967-:8])+$signed(-{in[5175-:8],2'b0})+$signed({in[5183-:8],1'b0})+$signed(sharing126)+$signed(-1);
assign weighted_sum[483] = $signed(-{in[5191-:8],2'b0})+$signed({in[5199-:8],1'b0})+$signed({in[5207-:8],1'b0})+$signed(in[5207-:8])+$signed(-{in[5415-:8],3'b0})+$signed(-{in[5423-:8],3'b0})+$signed({in[4975-:8],1'b0})+$signed({in[4983-:8],2'b0})+$signed(-{in[5431-:8],1'b0})+$signed(in[4983-:8])+$signed(sharing127)+$signed(-1);
assign weighted_sum[484] = $signed({in[4999-:8],2'b0})+$signed(-{in[5447-:8],1'b0})+$signed(in[4999-:8])+$signed(-{in[5207-:8],2'b0})+$signed({in[5215-:8],1'b0})+$signed({in[5223-:8],1'b0})+$signed(in[5223-:8])+$signed(-{in[5431-:8],3'b0})+$signed(-{in[5439-:8],3'b0})+$signed({in[4991-:8],1'b0})+$signed(sharing128)+$signed(-1);
assign weighted_sum[485] = $signed(-{in[5447-:8],3'b0})+$signed(-{in[5455-:8],3'b0})+$signed({in[5007-:8],1'b0})+$signed({in[5015-:8],2'b0})+$signed(-{in[5463-:8],1'b0})+$signed(in[5015-:8])+$signed(-{in[5223-:8],2'b0})+$signed({in[5231-:8],1'b0})+$signed({in[5239-:8],1'b0})+$signed(in[5239-:8])+$signed(sharing129)+$signed(-1);
assign weighted_sum[486] = $signed({in[5255-:8],1'b0})+$signed(in[5255-:8])+$signed(-{in[5463-:8],3'b0})+$signed(-{in[5471-:8],3'b0})+$signed({in[5023-:8],1'b0})+$signed({in[5031-:8],2'b0})+$signed(-{in[5479-:8],1'b0})+$signed(in[5031-:8])+$signed(-{in[5239-:8],2'b0})+$signed({in[5247-:8],1'b0})+$signed(sharing130)+$signed(-1);
assign weighted_sum[487] = $signed(-{in[5255-:8],2'b0})+$signed({in[5263-:8],1'b0})+$signed({in[5271-:8],1'b0})+$signed(in[5271-:8])+$signed(-{in[5479-:8],3'b0})+$signed(-{in[5487-:8],3'b0})+$signed({in[5039-:8],1'b0})+$signed({in[5047-:8],2'b0})+$signed(-{in[5495-:8],1'b0})+$signed(in[5047-:8])+$signed(sharing131)+$signed(-1);
assign weighted_sum[488] = $signed({in[5063-:8],2'b0})+$signed(-{in[5511-:8],1'b0})+$signed(in[5063-:8])+$signed(-{in[5271-:8],2'b0})+$signed({in[5279-:8],1'b0})+$signed({in[5287-:8],1'b0})+$signed(in[5287-:8])+$signed(-{in[5495-:8],3'b0})+$signed(-{in[5503-:8],3'b0})+$signed({in[5055-:8],1'b0})+$signed(sharing166)+$signed(-1);
assign weighted_sum[489] = $signed(-{in[5511-:8],3'b0})+$signed(-{in[5519-:8],3'b0})+$signed({in[5071-:8],1'b0})+$signed({in[5079-:8],2'b0})+$signed(-{in[5527-:8],1'b0})+$signed(in[5079-:8])+$signed(-{in[5287-:8],2'b0})+$signed({in[5295-:8],1'b0})+$signed({in[5303-:8],1'b0})+$signed(in[5303-:8])+$signed(sharing132)+$signed(-1);
assign weighted_sum[490] = $signed({in[5319-:8],1'b0})+$signed(in[5319-:8])+$signed(-{in[5527-:8],3'b0})+$signed(-{in[5535-:8],3'b0})+$signed({in[5087-:8],1'b0})+$signed({in[5095-:8],2'b0})+$signed(-{in[5543-:8],1'b0})+$signed(in[5095-:8])+$signed(-{in[5303-:8],2'b0})+$signed({in[5311-:8],1'b0})+$signed(sharing133)+$signed(-1);
assign weighted_sum[491] = $signed(-{in[5319-:8],2'b0})+$signed({in[5327-:8],1'b0})+$signed({in[5335-:8],1'b0})+$signed(in[5335-:8])+$signed(-{in[5543-:8],3'b0})+$signed(-{in[5551-:8],3'b0})+$signed({in[5103-:8],1'b0})+$signed({in[5111-:8],2'b0})+$signed(-{in[5559-:8],1'b0})+$signed(in[5111-:8])+$signed(sharing134)+$signed(-1);
assign weighted_sum[492] = $signed({in[5127-:8],2'b0})+$signed(-{in[5575-:8],1'b0})+$signed(in[5127-:8])+$signed(-{in[5335-:8],2'b0})+$signed({in[5343-:8],1'b0})+$signed({in[5351-:8],1'b0})+$signed(in[5351-:8])+$signed(-{in[5559-:8],3'b0})+$signed(-{in[5567-:8],3'b0})+$signed({in[5119-:8],1'b0})+$signed(sharing135)+$signed(-1);
assign weighted_sum[493] = $signed(-{in[5575-:8],3'b0})+$signed(-{in[5583-:8],3'b0})+$signed({in[5135-:8],1'b0})+$signed({in[5143-:8],2'b0})+$signed(-{in[5591-:8],1'b0})+$signed(in[5143-:8])+$signed(-{in[5351-:8],2'b0})+$signed({in[5359-:8],1'b0})+$signed({in[5367-:8],1'b0})+$signed(in[5367-:8])+$signed(sharing136)+$signed(-1);
assign weighted_sum[494] = $signed(-{in[5831-:8],3'b0})+$signed(-{in[5839-:8],3'b0})+$signed({in[5391-:8],1'b0})+$signed({in[5399-:8],2'b0})+$signed(-{in[5847-:8],1'b0})+$signed(in[5399-:8])+$signed(-{in[5607-:8],2'b0})+$signed({in[5615-:8],1'b0})+$signed({in[5623-:8],1'b0})+$signed(in[5623-:8])+$signed(sharing137)+$signed(-1);
assign weighted_sum[495] = $signed({in[5639-:8],1'b0})+$signed(in[5639-:8])+$signed(-{in[5847-:8],3'b0})+$signed(-{in[5855-:8],3'b0})+$signed({in[5407-:8],1'b0})+$signed({in[5415-:8],2'b0})+$signed(-{in[5863-:8],1'b0})+$signed(in[5415-:8])+$signed(-{in[5623-:8],2'b0})+$signed({in[5631-:8],1'b0})+$signed(sharing138)+$signed(-1);
assign weighted_sum[496] = $signed(-{in[5639-:8],2'b0})+$signed({in[5647-:8],1'b0})+$signed({in[5655-:8],1'b0})+$signed(in[5655-:8])+$signed(-{in[5863-:8],3'b0})+$signed(-{in[5871-:8],3'b0})+$signed({in[5423-:8],1'b0})+$signed({in[5431-:8],2'b0})+$signed(-{in[5879-:8],1'b0})+$signed(in[5431-:8])+$signed(sharing167)+$signed(-1);
assign weighted_sum[497] = $signed({in[5447-:8],2'b0})+$signed(-{in[5895-:8],1'b0})+$signed(in[5447-:8])+$signed(-{in[5655-:8],2'b0})+$signed({in[5663-:8],1'b0})+$signed({in[5671-:8],1'b0})+$signed(in[5671-:8])+$signed(-{in[5879-:8],3'b0})+$signed(-{in[5887-:8],3'b0})+$signed({in[5439-:8],1'b0})+$signed(sharing139)+$signed(-1);
assign weighted_sum[498] = $signed(-{in[5895-:8],3'b0})+$signed(-{in[5903-:8],3'b0})+$signed({in[5455-:8],1'b0})+$signed({in[5463-:8],2'b0})+$signed(-{in[5911-:8],1'b0})+$signed(in[5463-:8])+$signed(-{in[5671-:8],2'b0})+$signed({in[5679-:8],1'b0})+$signed({in[5687-:8],1'b0})+$signed(in[5687-:8])+$signed(sharing140)+$signed(-1);
assign weighted_sum[499] = $signed({in[5703-:8],1'b0})+$signed(in[5703-:8])+$signed(-{in[5911-:8],3'b0})+$signed(-{in[5919-:8],3'b0})+$signed({in[5471-:8],1'b0})+$signed({in[5479-:8],2'b0})+$signed(-{in[5927-:8],1'b0})+$signed(in[5479-:8])+$signed(-{in[5687-:8],2'b0})+$signed({in[5695-:8],1'b0})+$signed(sharing141)+$signed(-1);
assign weighted_sum[500] = $signed(-{in[5703-:8],2'b0})+$signed({in[5711-:8],1'b0})+$signed({in[5719-:8],1'b0})+$signed(in[5719-:8])+$signed(-{in[5927-:8],3'b0})+$signed(-{in[5935-:8],3'b0})+$signed({in[5487-:8],1'b0})+$signed({in[5495-:8],2'b0})+$signed(-{in[5943-:8],1'b0})+$signed(in[5495-:8])+$signed(sharing142)+$signed(-1);
assign weighted_sum[501] = $signed({in[5511-:8],2'b0})+$signed(-{in[5959-:8],1'b0})+$signed(in[5511-:8])+$signed(-{in[5719-:8],2'b0})+$signed({in[5727-:8],1'b0})+$signed({in[5735-:8],1'b0})+$signed(in[5735-:8])+$signed(-{in[5943-:8],3'b0})+$signed(-{in[5951-:8],3'b0})+$signed({in[5503-:8],1'b0})+$signed(sharing143)+$signed(-1);
assign weighted_sum[502] = $signed(-{in[5959-:8],3'b0})+$signed(-{in[5967-:8],3'b0})+$signed({in[5519-:8],1'b0})+$signed({in[5527-:8],2'b0})+$signed(-{in[5975-:8],1'b0})+$signed(in[5527-:8])+$signed(-{in[5735-:8],2'b0})+$signed({in[5743-:8],1'b0})+$signed({in[5751-:8],1'b0})+$signed(in[5751-:8])+$signed(sharing144)+$signed(-1);
assign weighted_sum[503] = $signed({in[5767-:8],1'b0})+$signed(in[5767-:8])+$signed(-{in[5975-:8],3'b0})+$signed(-{in[5983-:8],3'b0})+$signed({in[5535-:8],1'b0})+$signed({in[5543-:8],2'b0})+$signed(-{in[5991-:8],1'b0})+$signed(in[5543-:8])+$signed(-{in[5751-:8],2'b0})+$signed({in[5759-:8],1'b0})+$signed(sharing145)+$signed(-1);
assign weighted_sum[504] = $signed(-{in[5767-:8],2'b0})+$signed({in[5775-:8],1'b0})+$signed({in[5783-:8],1'b0})+$signed(in[5783-:8])+$signed(-{in[5991-:8],3'b0})+$signed(-{in[5999-:8],3'b0})+$signed({in[5551-:8],1'b0})+$signed({in[5559-:8],2'b0})+$signed(-{in[6007-:8],1'b0})+$signed(in[5559-:8])+$signed(sharing168)+$signed(-1);
assign weighted_sum[505] = $signed({in[5575-:8],2'b0})+$signed(-{in[6023-:8],1'b0})+$signed(in[5575-:8])+$signed(-{in[5783-:8],2'b0})+$signed({in[5791-:8],1'b0})+$signed({in[5799-:8],1'b0})+$signed(in[5799-:8])+$signed(-{in[6007-:8],3'b0})+$signed(-{in[6015-:8],3'b0})+$signed({in[5567-:8],1'b0})+$signed(sharing146)+$signed(-1);
assign weighted_sum[506] = $signed(-{in[6023-:8],3'b0})+$signed(-{in[6031-:8],3'b0})+$signed({in[5583-:8],1'b0})+$signed({in[5591-:8],2'b0})+$signed(-{in[6039-:8],1'b0})+$signed(in[5591-:8])+$signed(-{in[5799-:8],2'b0})+$signed({in[5807-:8],1'b0})+$signed({in[5815-:8],1'b0})+$signed(in[5815-:8])+$signed(sharing147)+$signed(-1);
assign relu_out[0] = (weighted_sum[0][12]==1) ? 4'd0 : (weighted_sum[0][11:8] > 6 ? 4'd6 : weighted_sum[0][11:8]);
assign relu_out[1] = (weighted_sum[1][12]==1) ? 4'd0 : (weighted_sum[1][11:8] > 6 ? 4'd6 : weighted_sum[1][11:8]);
assign relu_out[2] = (weighted_sum[2][12]==1) ? 4'd0 : (weighted_sum[2][11:8] > 6 ? 4'd6 : weighted_sum[2][11:8]);
assign relu_out[3] = (weighted_sum[3][12]==1) ? 4'd0 : (weighted_sum[3][11:8] > 6 ? 4'd6 : weighted_sum[3][11:8]);
assign relu_out[4] = (weighted_sum[4][12]==1) ? 4'd0 : (weighted_sum[4][11:8] > 6 ? 4'd6 : weighted_sum[4][11:8]);
assign relu_out[5] = (weighted_sum[5][12]==1) ? 4'd0 : (weighted_sum[5][11:8] > 6 ? 4'd6 : weighted_sum[5][11:8]);
assign relu_out[6] = (weighted_sum[6][12]==1) ? 4'd0 : (weighted_sum[6][11:8] > 6 ? 4'd6 : weighted_sum[6][11:8]);
assign relu_out[7] = (weighted_sum[7][12]==1) ? 4'd0 : (weighted_sum[7][11:8] > 6 ? 4'd6 : weighted_sum[7][11:8]);
assign relu_out[8] = (weighted_sum[8][12]==1) ? 4'd0 : (weighted_sum[8][11:8] > 6 ? 4'd6 : weighted_sum[8][11:8]);
assign relu_out[9] = (weighted_sum[9][12]==1) ? 4'd0 : (weighted_sum[9][11:8] > 6 ? 4'd6 : weighted_sum[9][11:8]);
assign relu_out[10] = (weighted_sum[10][12]==1) ? 4'd0 : (weighted_sum[10][11:8] > 6 ? 4'd6 : weighted_sum[10][11:8]);
assign relu_out[11] = (weighted_sum[11][12]==1) ? 4'd0 : (weighted_sum[11][11:8] > 6 ? 4'd6 : weighted_sum[11][11:8]);
assign relu_out[12] = (weighted_sum[12][12]==1) ? 4'd0 : (weighted_sum[12][11:8] > 6 ? 4'd6 : weighted_sum[12][11:8]);
assign relu_out[13] = (weighted_sum[13][12]==1) ? 4'd0 : (weighted_sum[13][11:8] > 6 ? 4'd6 : weighted_sum[13][11:8]);
assign relu_out[14] = (weighted_sum[14][12]==1) ? 4'd0 : (weighted_sum[14][11:8] > 6 ? 4'd6 : weighted_sum[14][11:8]);
assign relu_out[15] = (weighted_sum[15][12]==1) ? 4'd0 : (weighted_sum[15][11:8] > 6 ? 4'd6 : weighted_sum[15][11:8]);
assign relu_out[16] = (weighted_sum[16][12]==1) ? 4'd0 : (weighted_sum[16][11:8] > 6 ? 4'd6 : weighted_sum[16][11:8]);
assign relu_out[17] = (weighted_sum[17][12]==1) ? 4'd0 : (weighted_sum[17][11:8] > 6 ? 4'd6 : weighted_sum[17][11:8]);
assign relu_out[18] = (weighted_sum[18][12]==1) ? 4'd0 : (weighted_sum[18][11:8] > 6 ? 4'd6 : weighted_sum[18][11:8]);
assign relu_out[19] = (weighted_sum[19][12]==1) ? 4'd0 : (weighted_sum[19][11:8] > 6 ? 4'd6 : weighted_sum[19][11:8]);
assign relu_out[20] = (weighted_sum[20][12]==1) ? 4'd0 : (weighted_sum[20][11:8] > 6 ? 4'd6 : weighted_sum[20][11:8]);
assign relu_out[21] = (weighted_sum[21][12]==1) ? 4'd0 : (weighted_sum[21][11:8] > 6 ? 4'd6 : weighted_sum[21][11:8]);
assign relu_out[22] = (weighted_sum[22][12]==1) ? 4'd0 : (weighted_sum[22][11:8] > 6 ? 4'd6 : weighted_sum[22][11:8]);
assign relu_out[23] = (weighted_sum[23][12]==1) ? 4'd0 : (weighted_sum[23][11:8] > 6 ? 4'd6 : weighted_sum[23][11:8]);
assign relu_out[24] = (weighted_sum[24][12]==1) ? 4'd0 : (weighted_sum[24][11:8] > 6 ? 4'd6 : weighted_sum[24][11:8]);
assign relu_out[25] = (weighted_sum[25][12]==1) ? 4'd0 : (weighted_sum[25][11:8] > 6 ? 4'd6 : weighted_sum[25][11:8]);
assign relu_out[26] = (weighted_sum[26][12]==1) ? 4'd0 : (weighted_sum[26][11:8] > 6 ? 4'd6 : weighted_sum[26][11:8]);
assign relu_out[27] = (weighted_sum[27][12]==1) ? 4'd0 : (weighted_sum[27][11:8] > 6 ? 4'd6 : weighted_sum[27][11:8]);
assign relu_out[28] = (weighted_sum[28][12]==1) ? 4'd0 : (weighted_sum[28][11:8] > 6 ? 4'd6 : weighted_sum[28][11:8]);
assign relu_out[29] = (weighted_sum[29][12]==1) ? 4'd0 : (weighted_sum[29][11:8] > 6 ? 4'd6 : weighted_sum[29][11:8]);
assign relu_out[30] = (weighted_sum[30][12]==1) ? 4'd0 : (weighted_sum[30][11:8] > 6 ? 4'd6 : weighted_sum[30][11:8]);
assign relu_out[31] = (weighted_sum[31][12]==1) ? 4'd0 : (weighted_sum[31][11:8] > 6 ? 4'd6 : weighted_sum[31][11:8]);
assign relu_out[32] = (weighted_sum[32][12]==1) ? 4'd0 : (weighted_sum[32][11:8] > 6 ? 4'd6 : weighted_sum[32][11:8]);
assign relu_out[33] = (weighted_sum[33][12]==1) ? 4'd0 : (weighted_sum[33][11:8] > 6 ? 4'd6 : weighted_sum[33][11:8]);
assign relu_out[34] = (weighted_sum[34][12]==1) ? 4'd0 : (weighted_sum[34][11:8] > 6 ? 4'd6 : weighted_sum[34][11:8]);
assign relu_out[35] = (weighted_sum[35][12]==1) ? 4'd0 : (weighted_sum[35][11:8] > 6 ? 4'd6 : weighted_sum[35][11:8]);
assign relu_out[36] = (weighted_sum[36][12]==1) ? 4'd0 : (weighted_sum[36][11:8] > 6 ? 4'd6 : weighted_sum[36][11:8]);
assign relu_out[37] = (weighted_sum[37][12]==1) ? 4'd0 : (weighted_sum[37][11:8] > 6 ? 4'd6 : weighted_sum[37][11:8]);
assign relu_out[38] = (weighted_sum[38][12]==1) ? 4'd0 : (weighted_sum[38][11:8] > 6 ? 4'd6 : weighted_sum[38][11:8]);
assign relu_out[39] = (weighted_sum[39][12]==1) ? 4'd0 : (weighted_sum[39][11:8] > 6 ? 4'd6 : weighted_sum[39][11:8]);
assign relu_out[40] = (weighted_sum[40][12]==1) ? 4'd0 : (weighted_sum[40][11:8] > 6 ? 4'd6 : weighted_sum[40][11:8]);
assign relu_out[41] = (weighted_sum[41][12]==1) ? 4'd0 : (weighted_sum[41][11:8] > 6 ? 4'd6 : weighted_sum[41][11:8]);
assign relu_out[42] = (weighted_sum[42][12]==1) ? 4'd0 : (weighted_sum[42][11:8] > 6 ? 4'd6 : weighted_sum[42][11:8]);
assign relu_out[43] = (weighted_sum[43][12]==1) ? 4'd0 : (weighted_sum[43][11:8] > 6 ? 4'd6 : weighted_sum[43][11:8]);
assign relu_out[44] = (weighted_sum[44][12]==1) ? 4'd0 : (weighted_sum[44][11:8] > 6 ? 4'd6 : weighted_sum[44][11:8]);
assign relu_out[45] = (weighted_sum[45][12]==1) ? 4'd0 : (weighted_sum[45][11:8] > 6 ? 4'd6 : weighted_sum[45][11:8]);
assign relu_out[46] = (weighted_sum[46][12]==1) ? 4'd0 : (weighted_sum[46][11:8] > 6 ? 4'd6 : weighted_sum[46][11:8]);
assign relu_out[47] = (weighted_sum[47][12]==1) ? 4'd0 : (weighted_sum[47][11:8] > 6 ? 4'd6 : weighted_sum[47][11:8]);
assign relu_out[48] = (weighted_sum[48][12]==1) ? 4'd0 : (weighted_sum[48][11:8] > 6 ? 4'd6 : weighted_sum[48][11:8]);
assign relu_out[49] = (weighted_sum[49][12]==1) ? 4'd0 : (weighted_sum[49][11:8] > 6 ? 4'd6 : weighted_sum[49][11:8]);
assign relu_out[50] = (weighted_sum[50][12]==1) ? 4'd0 : (weighted_sum[50][11:8] > 6 ? 4'd6 : weighted_sum[50][11:8]);
assign relu_out[51] = (weighted_sum[51][12]==1) ? 4'd0 : (weighted_sum[51][11:8] > 6 ? 4'd6 : weighted_sum[51][11:8]);
assign relu_out[52] = (weighted_sum[52][12]==1) ? 4'd0 : (weighted_sum[52][11:8] > 6 ? 4'd6 : weighted_sum[52][11:8]);
assign relu_out[53] = (weighted_sum[53][12]==1) ? 4'd0 : (weighted_sum[53][11:8] > 6 ? 4'd6 : weighted_sum[53][11:8]);
assign relu_out[54] = (weighted_sum[54][12]==1) ? 4'd0 : (weighted_sum[54][11:8] > 6 ? 4'd6 : weighted_sum[54][11:8]);
assign relu_out[55] = (weighted_sum[55][12]==1) ? 4'd0 : (weighted_sum[55][11:8] > 6 ? 4'd6 : weighted_sum[55][11:8]);
assign relu_out[56] = (weighted_sum[56][12]==1) ? 4'd0 : (weighted_sum[56][11:8] > 6 ? 4'd6 : weighted_sum[56][11:8]);
assign relu_out[57] = (weighted_sum[57][12]==1) ? 4'd0 : (weighted_sum[57][11:8] > 6 ? 4'd6 : weighted_sum[57][11:8]);
assign relu_out[58] = (weighted_sum[58][12]==1) ? 4'd0 : (weighted_sum[58][11:8] > 6 ? 4'd6 : weighted_sum[58][11:8]);
assign relu_out[59] = (weighted_sum[59][12]==1) ? 4'd0 : (weighted_sum[59][11:8] > 6 ? 4'd6 : weighted_sum[59][11:8]);
assign relu_out[60] = (weighted_sum[60][12]==1) ? 4'd0 : (weighted_sum[60][11:8] > 6 ? 4'd6 : weighted_sum[60][11:8]);
assign relu_out[61] = (weighted_sum[61][12]==1) ? 4'd0 : (weighted_sum[61][11:8] > 6 ? 4'd6 : weighted_sum[61][11:8]);
assign relu_out[62] = (weighted_sum[62][12]==1) ? 4'd0 : (weighted_sum[62][11:8] > 6 ? 4'd6 : weighted_sum[62][11:8]);
assign relu_out[63] = (weighted_sum[63][12]==1) ? 4'd0 : (weighted_sum[63][11:8] > 6 ? 4'd6 : weighted_sum[63][11:8]);
assign relu_out[64] = (weighted_sum[64][12]==1) ? 4'd0 : (weighted_sum[64][11:8] > 6 ? 4'd6 : weighted_sum[64][11:8]);
assign relu_out[65] = (weighted_sum[65][12]==1) ? 4'd0 : (weighted_sum[65][11:8] > 6 ? 4'd6 : weighted_sum[65][11:8]);
assign relu_out[66] = (weighted_sum[66][12]==1) ? 4'd0 : (weighted_sum[66][11:8] > 6 ? 4'd6 : weighted_sum[66][11:8]);
assign relu_out[67] = (weighted_sum[67][12]==1) ? 4'd0 : (weighted_sum[67][11:8] > 6 ? 4'd6 : weighted_sum[67][11:8]);
assign relu_out[68] = (weighted_sum[68][12]==1) ? 4'd0 : (weighted_sum[68][11:8] > 6 ? 4'd6 : weighted_sum[68][11:8]);
assign relu_out[69] = (weighted_sum[69][12]==1) ? 4'd0 : (weighted_sum[69][11:8] > 6 ? 4'd6 : weighted_sum[69][11:8]);
assign relu_out[70] = (weighted_sum[70][12]==1) ? 4'd0 : (weighted_sum[70][11:8] > 6 ? 4'd6 : weighted_sum[70][11:8]);
assign relu_out[71] = (weighted_sum[71][12]==1) ? 4'd0 : (weighted_sum[71][11:8] > 6 ? 4'd6 : weighted_sum[71][11:8]);
assign relu_out[72] = (weighted_sum[72][12]==1) ? 4'd0 : (weighted_sum[72][11:8] > 6 ? 4'd6 : weighted_sum[72][11:8]);
assign relu_out[73] = (weighted_sum[73][12]==1) ? 4'd0 : (weighted_sum[73][11:8] > 6 ? 4'd6 : weighted_sum[73][11:8]);
assign relu_out[74] = (weighted_sum[74][12]==1) ? 4'd0 : (weighted_sum[74][11:8] > 6 ? 4'd6 : weighted_sum[74][11:8]);
assign relu_out[75] = (weighted_sum[75][12]==1) ? 4'd0 : (weighted_sum[75][11:8] > 6 ? 4'd6 : weighted_sum[75][11:8]);
assign relu_out[76] = (weighted_sum[76][12]==1) ? 4'd0 : (weighted_sum[76][11:8] > 6 ? 4'd6 : weighted_sum[76][11:8]);
assign relu_out[77] = (weighted_sum[77][12]==1) ? 4'd0 : (weighted_sum[77][11:8] > 6 ? 4'd6 : weighted_sum[77][11:8]);
assign relu_out[78] = (weighted_sum[78][12]==1) ? 4'd0 : (weighted_sum[78][11:8] > 6 ? 4'd6 : weighted_sum[78][11:8]);
assign relu_out[79] = (weighted_sum[79][12]==1) ? 4'd0 : (weighted_sum[79][11:8] > 6 ? 4'd6 : weighted_sum[79][11:8]);
assign relu_out[80] = (weighted_sum[80][12]==1) ? 4'd0 : (weighted_sum[80][11:8] > 6 ? 4'd6 : weighted_sum[80][11:8]);
assign relu_out[81] = (weighted_sum[81][12]==1) ? 4'd0 : (weighted_sum[81][11:8] > 6 ? 4'd6 : weighted_sum[81][11:8]);
assign relu_out[82] = (weighted_sum[82][12]==1) ? 4'd0 : (weighted_sum[82][11:8] > 6 ? 4'd6 : weighted_sum[82][11:8]);
assign relu_out[83] = (weighted_sum[83][12]==1) ? 4'd0 : (weighted_sum[83][11:8] > 6 ? 4'd6 : weighted_sum[83][11:8]);
assign relu_out[84] = (weighted_sum[84][12]==1) ? 4'd0 : (weighted_sum[84][11:8] > 6 ? 4'd6 : weighted_sum[84][11:8]);
assign relu_out[85] = (weighted_sum[85][12]==1) ? 4'd0 : (weighted_sum[85][11:8] > 6 ? 4'd6 : weighted_sum[85][11:8]);
assign relu_out[86] = (weighted_sum[86][12]==1) ? 4'd0 : (weighted_sum[86][11:8] > 6 ? 4'd6 : weighted_sum[86][11:8]);
assign relu_out[87] = (weighted_sum[87][12]==1) ? 4'd0 : (weighted_sum[87][11:8] > 6 ? 4'd6 : weighted_sum[87][11:8]);
assign relu_out[88] = (weighted_sum[88][12]==1) ? 4'd0 : (weighted_sum[88][11:8] > 6 ? 4'd6 : weighted_sum[88][11:8]);
assign relu_out[89] = (weighted_sum[89][12]==1) ? 4'd0 : (weighted_sum[89][11:8] > 6 ? 4'd6 : weighted_sum[89][11:8]);
assign relu_out[90] = (weighted_sum[90][12]==1) ? 4'd0 : (weighted_sum[90][11:8] > 6 ? 4'd6 : weighted_sum[90][11:8]);
assign relu_out[91] = (weighted_sum[91][12]==1) ? 4'd0 : (weighted_sum[91][11:8] > 6 ? 4'd6 : weighted_sum[91][11:8]);
assign relu_out[92] = (weighted_sum[92][12]==1) ? 4'd0 : (weighted_sum[92][11:8] > 6 ? 4'd6 : weighted_sum[92][11:8]);
assign relu_out[93] = (weighted_sum[93][12]==1) ? 4'd0 : (weighted_sum[93][11:8] > 6 ? 4'd6 : weighted_sum[93][11:8]);
assign relu_out[94] = (weighted_sum[94][12]==1) ? 4'd0 : (weighted_sum[94][11:8] > 6 ? 4'd6 : weighted_sum[94][11:8]);
assign relu_out[95] = (weighted_sum[95][12]==1) ? 4'd0 : (weighted_sum[95][11:8] > 6 ? 4'd6 : weighted_sum[95][11:8]);
assign relu_out[96] = (weighted_sum[96][12]==1) ? 4'd0 : (weighted_sum[96][11:8] > 6 ? 4'd6 : weighted_sum[96][11:8]);
assign relu_out[97] = (weighted_sum[97][12]==1) ? 4'd0 : (weighted_sum[97][11:8] > 6 ? 4'd6 : weighted_sum[97][11:8]);
assign relu_out[98] = (weighted_sum[98][12]==1) ? 4'd0 : (weighted_sum[98][11:8] > 6 ? 4'd6 : weighted_sum[98][11:8]);
assign relu_out[99] = (weighted_sum[99][12]==1) ? 4'd0 : (weighted_sum[99][11:8] > 6 ? 4'd6 : weighted_sum[99][11:8]);
assign relu_out[100] = (weighted_sum[100][12]==1) ? 4'd0 : (weighted_sum[100][11:8] > 6 ? 4'd6 : weighted_sum[100][11:8]);
assign relu_out[101] = (weighted_sum[101][12]==1) ? 4'd0 : (weighted_sum[101][11:8] > 6 ? 4'd6 : weighted_sum[101][11:8]);
assign relu_out[102] = (weighted_sum[102][12]==1) ? 4'd0 : (weighted_sum[102][11:8] > 6 ? 4'd6 : weighted_sum[102][11:8]);
assign relu_out[103] = (weighted_sum[103][12]==1) ? 4'd0 : (weighted_sum[103][11:8] > 6 ? 4'd6 : weighted_sum[103][11:8]);
assign relu_out[104] = (weighted_sum[104][12]==1) ? 4'd0 : (weighted_sum[104][11:8] > 6 ? 4'd6 : weighted_sum[104][11:8]);
assign relu_out[105] = (weighted_sum[105][12]==1) ? 4'd0 : (weighted_sum[105][11:8] > 6 ? 4'd6 : weighted_sum[105][11:8]);
assign relu_out[106] = (weighted_sum[106][12]==1) ? 4'd0 : (weighted_sum[106][11:8] > 6 ? 4'd6 : weighted_sum[106][11:8]);
assign relu_out[107] = (weighted_sum[107][12]==1) ? 4'd0 : (weighted_sum[107][11:8] > 6 ? 4'd6 : weighted_sum[107][11:8]);
assign relu_out[108] = (weighted_sum[108][12]==1) ? 4'd0 : (weighted_sum[108][11:8] > 6 ? 4'd6 : weighted_sum[108][11:8]);
assign relu_out[109] = (weighted_sum[109][12]==1) ? 4'd0 : (weighted_sum[109][11:8] > 6 ? 4'd6 : weighted_sum[109][11:8]);
assign relu_out[110] = (weighted_sum[110][12]==1) ? 4'd0 : (weighted_sum[110][11:8] > 6 ? 4'd6 : weighted_sum[110][11:8]);
assign relu_out[111] = (weighted_sum[111][12]==1) ? 4'd0 : (weighted_sum[111][11:8] > 6 ? 4'd6 : weighted_sum[111][11:8]);
assign relu_out[112] = (weighted_sum[112][12]==1) ? 4'd0 : (weighted_sum[112][11:8] > 6 ? 4'd6 : weighted_sum[112][11:8]);
assign relu_out[113] = (weighted_sum[113][12]==1) ? 4'd0 : (weighted_sum[113][11:8] > 6 ? 4'd6 : weighted_sum[113][11:8]);
assign relu_out[114] = (weighted_sum[114][12]==1) ? 4'd0 : (weighted_sum[114][11:8] > 6 ? 4'd6 : weighted_sum[114][11:8]);
assign relu_out[115] = (weighted_sum[115][12]==1) ? 4'd0 : (weighted_sum[115][11:8] > 6 ? 4'd6 : weighted_sum[115][11:8]);
assign relu_out[116] = (weighted_sum[116][12]==1) ? 4'd0 : (weighted_sum[116][11:8] > 6 ? 4'd6 : weighted_sum[116][11:8]);
assign relu_out[117] = (weighted_sum[117][12]==1) ? 4'd0 : (weighted_sum[117][11:8] > 6 ? 4'd6 : weighted_sum[117][11:8]);
assign relu_out[118] = (weighted_sum[118][12]==1) ? 4'd0 : (weighted_sum[118][11:8] > 6 ? 4'd6 : weighted_sum[118][11:8]);
assign relu_out[119] = (weighted_sum[119][12]==1) ? 4'd0 : (weighted_sum[119][11:8] > 6 ? 4'd6 : weighted_sum[119][11:8]);
assign relu_out[120] = (weighted_sum[120][12]==1) ? 4'd0 : (weighted_sum[120][11:8] > 6 ? 4'd6 : weighted_sum[120][11:8]);
assign relu_out[121] = (weighted_sum[121][12]==1) ? 4'd0 : (weighted_sum[121][11:8] > 6 ? 4'd6 : weighted_sum[121][11:8]);
assign relu_out[122] = (weighted_sum[122][12]==1) ? 4'd0 : (weighted_sum[122][11:8] > 6 ? 4'd6 : weighted_sum[122][11:8]);
assign relu_out[123] = (weighted_sum[123][12]==1) ? 4'd0 : (weighted_sum[123][11:8] > 6 ? 4'd6 : weighted_sum[123][11:8]);
assign relu_out[124] = (weighted_sum[124][12]==1) ? 4'd0 : (weighted_sum[124][11:8] > 6 ? 4'd6 : weighted_sum[124][11:8]);
assign relu_out[125] = (weighted_sum[125][12]==1) ? 4'd0 : (weighted_sum[125][11:8] > 6 ? 4'd6 : weighted_sum[125][11:8]);
assign relu_out[126] = (weighted_sum[126][12]==1) ? 4'd0 : (weighted_sum[126][11:8] > 6 ? 4'd6 : weighted_sum[126][11:8]);
assign relu_out[127] = (weighted_sum[127][12]==1) ? 4'd0 : (weighted_sum[127][11:8] > 6 ? 4'd6 : weighted_sum[127][11:8]);
assign relu_out[128] = (weighted_sum[128][12]==1) ? 4'd0 : (weighted_sum[128][11:8] > 6 ? 4'd6 : weighted_sum[128][11:8]);
assign relu_out[129] = (weighted_sum[129][12]==1) ? 4'd0 : (weighted_sum[129][11:8] > 6 ? 4'd6 : weighted_sum[129][11:8]);
assign relu_out[130] = (weighted_sum[130][12]==1) ? 4'd0 : (weighted_sum[130][11:8] > 6 ? 4'd6 : weighted_sum[130][11:8]);
assign relu_out[131] = (weighted_sum[131][12]==1) ? 4'd0 : (weighted_sum[131][11:8] > 6 ? 4'd6 : weighted_sum[131][11:8]);
assign relu_out[132] = (weighted_sum[132][12]==1) ? 4'd0 : (weighted_sum[132][11:8] > 6 ? 4'd6 : weighted_sum[132][11:8]);
assign relu_out[133] = (weighted_sum[133][12]==1) ? 4'd0 : (weighted_sum[133][11:8] > 6 ? 4'd6 : weighted_sum[133][11:8]);
assign relu_out[134] = (weighted_sum[134][12]==1) ? 4'd0 : (weighted_sum[134][11:8] > 6 ? 4'd6 : weighted_sum[134][11:8]);
assign relu_out[135] = (weighted_sum[135][12]==1) ? 4'd0 : (weighted_sum[135][11:8] > 6 ? 4'd6 : weighted_sum[135][11:8]);
assign relu_out[136] = (weighted_sum[136][12]==1) ? 4'd0 : (weighted_sum[136][11:8] > 6 ? 4'd6 : weighted_sum[136][11:8]);
assign relu_out[137] = (weighted_sum[137][12]==1) ? 4'd0 : (weighted_sum[137][11:8] > 6 ? 4'd6 : weighted_sum[137][11:8]);
assign relu_out[138] = (weighted_sum[138][12]==1) ? 4'd0 : (weighted_sum[138][11:8] > 6 ? 4'd6 : weighted_sum[138][11:8]);
assign relu_out[139] = (weighted_sum[139][12]==1) ? 4'd0 : (weighted_sum[139][11:8] > 6 ? 4'd6 : weighted_sum[139][11:8]);
assign relu_out[140] = (weighted_sum[140][12]==1) ? 4'd0 : (weighted_sum[140][11:8] > 6 ? 4'd6 : weighted_sum[140][11:8]);
assign relu_out[141] = (weighted_sum[141][12]==1) ? 4'd0 : (weighted_sum[141][11:8] > 6 ? 4'd6 : weighted_sum[141][11:8]);
assign relu_out[142] = (weighted_sum[142][12]==1) ? 4'd0 : (weighted_sum[142][11:8] > 6 ? 4'd6 : weighted_sum[142][11:8]);
assign relu_out[143] = (weighted_sum[143][12]==1) ? 4'd0 : (weighted_sum[143][11:8] > 6 ? 4'd6 : weighted_sum[143][11:8]);
assign relu_out[144] = (weighted_sum[144][12]==1) ? 4'd0 : (weighted_sum[144][11:8] > 6 ? 4'd6 : weighted_sum[144][11:8]);
assign relu_out[145] = (weighted_sum[145][12]==1) ? 4'd0 : (weighted_sum[145][11:8] > 6 ? 4'd6 : weighted_sum[145][11:8]);
assign relu_out[146] = (weighted_sum[146][12]==1) ? 4'd0 : (weighted_sum[146][11:8] > 6 ? 4'd6 : weighted_sum[146][11:8]);
assign relu_out[147] = (weighted_sum[147][12]==1) ? 4'd0 : (weighted_sum[147][11:8] > 6 ? 4'd6 : weighted_sum[147][11:8]);
assign relu_out[148] = (weighted_sum[148][12]==1) ? 4'd0 : (weighted_sum[148][11:8] > 6 ? 4'd6 : weighted_sum[148][11:8]);
assign relu_out[149] = (weighted_sum[149][12]==1) ? 4'd0 : (weighted_sum[149][11:8] > 6 ? 4'd6 : weighted_sum[149][11:8]);
assign relu_out[150] = (weighted_sum[150][12]==1) ? 4'd0 : (weighted_sum[150][11:8] > 6 ? 4'd6 : weighted_sum[150][11:8]);
assign relu_out[151] = (weighted_sum[151][12]==1) ? 4'd0 : (weighted_sum[151][11:8] > 6 ? 4'd6 : weighted_sum[151][11:8]);
assign relu_out[152] = (weighted_sum[152][12]==1) ? 4'd0 : (weighted_sum[152][11:8] > 6 ? 4'd6 : weighted_sum[152][11:8]);
assign relu_out[153] = (weighted_sum[153][12]==1) ? 4'd0 : (weighted_sum[153][11:8] > 6 ? 4'd6 : weighted_sum[153][11:8]);
assign relu_out[154] = (weighted_sum[154][12]==1) ? 4'd0 : (weighted_sum[154][11:8] > 6 ? 4'd6 : weighted_sum[154][11:8]);
assign relu_out[155] = (weighted_sum[155][12]==1) ? 4'd0 : (weighted_sum[155][11:8] > 6 ? 4'd6 : weighted_sum[155][11:8]);
assign relu_out[156] = (weighted_sum[156][12]==1) ? 4'd0 : (weighted_sum[156][11:8] > 6 ? 4'd6 : weighted_sum[156][11:8]);
assign relu_out[157] = (weighted_sum[157][12]==1) ? 4'd0 : (weighted_sum[157][11:8] > 6 ? 4'd6 : weighted_sum[157][11:8]);
assign relu_out[158] = (weighted_sum[158][12]==1) ? 4'd0 : (weighted_sum[158][11:8] > 6 ? 4'd6 : weighted_sum[158][11:8]);
assign relu_out[159] = (weighted_sum[159][12]==1) ? 4'd0 : (weighted_sum[159][11:8] > 6 ? 4'd6 : weighted_sum[159][11:8]);
assign relu_out[160] = (weighted_sum[160][12]==1) ? 4'd0 : (weighted_sum[160][11:8] > 6 ? 4'd6 : weighted_sum[160][11:8]);
assign relu_out[161] = (weighted_sum[161][12]==1) ? 4'd0 : (weighted_sum[161][11:8] > 6 ? 4'd6 : weighted_sum[161][11:8]);
assign relu_out[162] = (weighted_sum[162][12]==1) ? 4'd0 : (weighted_sum[162][11:8] > 6 ? 4'd6 : weighted_sum[162][11:8]);
assign relu_out[163] = (weighted_sum[163][12]==1) ? 4'd0 : (weighted_sum[163][11:8] > 6 ? 4'd6 : weighted_sum[163][11:8]);
assign relu_out[164] = (weighted_sum[164][12]==1) ? 4'd0 : (weighted_sum[164][11:8] > 6 ? 4'd6 : weighted_sum[164][11:8]);
assign relu_out[165] = (weighted_sum[165][12]==1) ? 4'd0 : (weighted_sum[165][11:8] > 6 ? 4'd6 : weighted_sum[165][11:8]);
assign relu_out[166] = (weighted_sum[166][12]==1) ? 4'd0 : (weighted_sum[166][11:8] > 6 ? 4'd6 : weighted_sum[166][11:8]);
assign relu_out[167] = (weighted_sum[167][12]==1) ? 4'd0 : (weighted_sum[167][11:8] > 6 ? 4'd6 : weighted_sum[167][11:8]);
assign relu_out[168] = (weighted_sum[168][12]==1) ? 4'd0 : (weighted_sum[168][11:8] > 6 ? 4'd6 : weighted_sum[168][11:8]);
assign relu_out[169] = (weighted_sum[169][12]==1) ? 4'd0 : (weighted_sum[169][11:8] > 6 ? 4'd6 : weighted_sum[169][11:8]);
assign relu_out[170] = (weighted_sum[170][12]==1) ? 4'd0 : (weighted_sum[170][11:8] > 6 ? 4'd6 : weighted_sum[170][11:8]);
assign relu_out[171] = (weighted_sum[171][12]==1) ? 4'd0 : (weighted_sum[171][11:8] > 6 ? 4'd6 : weighted_sum[171][11:8]);
assign relu_out[172] = (weighted_sum[172][12]==1) ? 4'd0 : (weighted_sum[172][11:8] > 6 ? 4'd6 : weighted_sum[172][11:8]);
assign relu_out[173] = (weighted_sum[173][12]==1) ? 4'd0 : (weighted_sum[173][11:8] > 6 ? 4'd6 : weighted_sum[173][11:8]);
assign relu_out[174] = (weighted_sum[174][12]==1) ? 4'd0 : (weighted_sum[174][11:8] > 6 ? 4'd6 : weighted_sum[174][11:8]);
assign relu_out[175] = (weighted_sum[175][12]==1) ? 4'd0 : (weighted_sum[175][11:8] > 6 ? 4'd6 : weighted_sum[175][11:8]);
assign relu_out[176] = (weighted_sum[176][12]==1) ? 4'd0 : (weighted_sum[176][11:8] > 6 ? 4'd6 : weighted_sum[176][11:8]);
assign relu_out[177] = (weighted_sum[177][12]==1) ? 4'd0 : (weighted_sum[177][11:8] > 6 ? 4'd6 : weighted_sum[177][11:8]);
assign relu_out[178] = (weighted_sum[178][12]==1) ? 4'd0 : (weighted_sum[178][11:8] > 6 ? 4'd6 : weighted_sum[178][11:8]);
assign relu_out[179] = (weighted_sum[179][12]==1) ? 4'd0 : (weighted_sum[179][11:8] > 6 ? 4'd6 : weighted_sum[179][11:8]);
assign relu_out[180] = (weighted_sum[180][12]==1) ? 4'd0 : (weighted_sum[180][11:8] > 6 ? 4'd6 : weighted_sum[180][11:8]);
assign relu_out[181] = (weighted_sum[181][12]==1) ? 4'd0 : (weighted_sum[181][11:8] > 6 ? 4'd6 : weighted_sum[181][11:8]);
assign relu_out[182] = (weighted_sum[182][12]==1) ? 4'd0 : (weighted_sum[182][11:8] > 6 ? 4'd6 : weighted_sum[182][11:8]);
assign relu_out[183] = (weighted_sum[183][12]==1) ? 4'd0 : (weighted_sum[183][11:8] > 6 ? 4'd6 : weighted_sum[183][11:8]);
assign relu_out[184] = (weighted_sum[184][12]==1) ? 4'd0 : (weighted_sum[184][11:8] > 6 ? 4'd6 : weighted_sum[184][11:8]);
assign relu_out[185] = (weighted_sum[185][12]==1) ? 4'd0 : (weighted_sum[185][11:8] > 6 ? 4'd6 : weighted_sum[185][11:8]);
assign relu_out[186] = (weighted_sum[186][12]==1) ? 4'd0 : (weighted_sum[186][11:8] > 6 ? 4'd6 : weighted_sum[186][11:8]);
assign relu_out[187] = (weighted_sum[187][12]==1) ? 4'd0 : (weighted_sum[187][11:8] > 6 ? 4'd6 : weighted_sum[187][11:8]);
assign relu_out[188] = (weighted_sum[188][12]==1) ? 4'd0 : (weighted_sum[188][11:8] > 6 ? 4'd6 : weighted_sum[188][11:8]);
assign relu_out[189] = (weighted_sum[189][12]==1) ? 4'd0 : (weighted_sum[189][11:8] > 6 ? 4'd6 : weighted_sum[189][11:8]);
assign relu_out[190] = (weighted_sum[190][12]==1) ? 4'd0 : (weighted_sum[190][11:8] > 6 ? 4'd6 : weighted_sum[190][11:8]);
assign relu_out[191] = (weighted_sum[191][12]==1) ? 4'd0 : (weighted_sum[191][11:8] > 6 ? 4'd6 : weighted_sum[191][11:8]);
assign relu_out[192] = (weighted_sum[192][12]==1) ? 4'd0 : (weighted_sum[192][11:8] > 6 ? 4'd6 : weighted_sum[192][11:8]);
assign relu_out[193] = (weighted_sum[193][12]==1) ? 4'd0 : (weighted_sum[193][11:8] > 6 ? 4'd6 : weighted_sum[193][11:8]);
assign relu_out[194] = (weighted_sum[194][12]==1) ? 4'd0 : (weighted_sum[194][11:8] > 6 ? 4'd6 : weighted_sum[194][11:8]);
assign relu_out[195] = (weighted_sum[195][12]==1) ? 4'd0 : (weighted_sum[195][11:8] > 6 ? 4'd6 : weighted_sum[195][11:8]);
assign relu_out[196] = (weighted_sum[196][12]==1) ? 4'd0 : (weighted_sum[196][11:8] > 6 ? 4'd6 : weighted_sum[196][11:8]);
assign relu_out[197] = (weighted_sum[197][12]==1) ? 4'd0 : (weighted_sum[197][11:8] > 6 ? 4'd6 : weighted_sum[197][11:8]);
assign relu_out[198] = (weighted_sum[198][12]==1) ? 4'd0 : (weighted_sum[198][11:8] > 6 ? 4'd6 : weighted_sum[198][11:8]);
assign relu_out[199] = (weighted_sum[199][12]==1) ? 4'd0 : (weighted_sum[199][11:8] > 6 ? 4'd6 : weighted_sum[199][11:8]);
assign relu_out[200] = (weighted_sum[200][12]==1) ? 4'd0 : (weighted_sum[200][11:8] > 6 ? 4'd6 : weighted_sum[200][11:8]);
assign relu_out[201] = (weighted_sum[201][12]==1) ? 4'd0 : (weighted_sum[201][11:8] > 6 ? 4'd6 : weighted_sum[201][11:8]);
assign relu_out[202] = (weighted_sum[202][12]==1) ? 4'd0 : (weighted_sum[202][11:8] > 6 ? 4'd6 : weighted_sum[202][11:8]);
assign relu_out[203] = (weighted_sum[203][12]==1) ? 4'd0 : (weighted_sum[203][11:8] > 6 ? 4'd6 : weighted_sum[203][11:8]);
assign relu_out[204] = (weighted_sum[204][12]==1) ? 4'd0 : (weighted_sum[204][11:8] > 6 ? 4'd6 : weighted_sum[204][11:8]);
assign relu_out[205] = (weighted_sum[205][12]==1) ? 4'd0 : (weighted_sum[205][11:8] > 6 ? 4'd6 : weighted_sum[205][11:8]);
assign relu_out[206] = (weighted_sum[206][12]==1) ? 4'd0 : (weighted_sum[206][11:8] > 6 ? 4'd6 : weighted_sum[206][11:8]);
assign relu_out[207] = (weighted_sum[207][12]==1) ? 4'd0 : (weighted_sum[207][11:8] > 6 ? 4'd6 : weighted_sum[207][11:8]);
assign relu_out[208] = (weighted_sum[208][12]==1) ? 4'd0 : (weighted_sum[208][11:8] > 6 ? 4'd6 : weighted_sum[208][11:8]);
assign relu_out[209] = (weighted_sum[209][12]==1) ? 4'd0 : (weighted_sum[209][11:8] > 6 ? 4'd6 : weighted_sum[209][11:8]);
assign relu_out[210] = (weighted_sum[210][12]==1) ? 4'd0 : (weighted_sum[210][11:8] > 6 ? 4'd6 : weighted_sum[210][11:8]);
assign relu_out[211] = (weighted_sum[211][12]==1) ? 4'd0 : (weighted_sum[211][11:8] > 6 ? 4'd6 : weighted_sum[211][11:8]);
assign relu_out[212] = (weighted_sum[212][12]==1) ? 4'd0 : (weighted_sum[212][11:8] > 6 ? 4'd6 : weighted_sum[212][11:8]);
assign relu_out[213] = (weighted_sum[213][12]==1) ? 4'd0 : (weighted_sum[213][11:8] > 6 ? 4'd6 : weighted_sum[213][11:8]);
assign relu_out[214] = (weighted_sum[214][12]==1) ? 4'd0 : (weighted_sum[214][11:8] > 6 ? 4'd6 : weighted_sum[214][11:8]);
assign relu_out[215] = (weighted_sum[215][12]==1) ? 4'd0 : (weighted_sum[215][11:8] > 6 ? 4'd6 : weighted_sum[215][11:8]);
assign relu_out[216] = (weighted_sum[216][12]==1) ? 4'd0 : (weighted_sum[216][11:8] > 6 ? 4'd6 : weighted_sum[216][11:8]);
assign relu_out[217] = (weighted_sum[217][12]==1) ? 4'd0 : (weighted_sum[217][11:8] > 6 ? 4'd6 : weighted_sum[217][11:8]);
assign relu_out[218] = (weighted_sum[218][12]==1) ? 4'd0 : (weighted_sum[218][11:8] > 6 ? 4'd6 : weighted_sum[218][11:8]);
assign relu_out[219] = (weighted_sum[219][12]==1) ? 4'd0 : (weighted_sum[219][11:8] > 6 ? 4'd6 : weighted_sum[219][11:8]);
assign relu_out[220] = (weighted_sum[220][12]==1) ? 4'd0 : (weighted_sum[220][11:8] > 6 ? 4'd6 : weighted_sum[220][11:8]);
assign relu_out[221] = (weighted_sum[221][12]==1) ? 4'd0 : (weighted_sum[221][11:8] > 6 ? 4'd6 : weighted_sum[221][11:8]);
assign relu_out[222] = (weighted_sum[222][12]==1) ? 4'd0 : (weighted_sum[222][11:8] > 6 ? 4'd6 : weighted_sum[222][11:8]);
assign relu_out[223] = (weighted_sum[223][12]==1) ? 4'd0 : (weighted_sum[223][11:8] > 6 ? 4'd6 : weighted_sum[223][11:8]);
assign relu_out[224] = (weighted_sum[224][12]==1) ? 4'd0 : (weighted_sum[224][11:8] > 6 ? 4'd6 : weighted_sum[224][11:8]);
assign relu_out[225] = (weighted_sum[225][12]==1) ? 4'd0 : (weighted_sum[225][11:8] > 6 ? 4'd6 : weighted_sum[225][11:8]);
assign relu_out[226] = (weighted_sum[226][12]==1) ? 4'd0 : (weighted_sum[226][11:8] > 6 ? 4'd6 : weighted_sum[226][11:8]);
assign relu_out[227] = (weighted_sum[227][12]==1) ? 4'd0 : (weighted_sum[227][11:8] > 6 ? 4'd6 : weighted_sum[227][11:8]);
assign relu_out[228] = (weighted_sum[228][12]==1) ? 4'd0 : (weighted_sum[228][11:8] > 6 ? 4'd6 : weighted_sum[228][11:8]);
assign relu_out[229] = (weighted_sum[229][12]==1) ? 4'd0 : (weighted_sum[229][11:8] > 6 ? 4'd6 : weighted_sum[229][11:8]);
assign relu_out[230] = (weighted_sum[230][12]==1) ? 4'd0 : (weighted_sum[230][11:8] > 6 ? 4'd6 : weighted_sum[230][11:8]);
assign relu_out[231] = (weighted_sum[231][12]==1) ? 4'd0 : (weighted_sum[231][11:8] > 6 ? 4'd6 : weighted_sum[231][11:8]);
assign relu_out[232] = (weighted_sum[232][12]==1) ? 4'd0 : (weighted_sum[232][11:8] > 6 ? 4'd6 : weighted_sum[232][11:8]);
assign relu_out[233] = (weighted_sum[233][12]==1) ? 4'd0 : (weighted_sum[233][11:8] > 6 ? 4'd6 : weighted_sum[233][11:8]);
assign relu_out[234] = (weighted_sum[234][12]==1) ? 4'd0 : (weighted_sum[234][11:8] > 6 ? 4'd6 : weighted_sum[234][11:8]);
assign relu_out[235] = (weighted_sum[235][12]==1) ? 4'd0 : (weighted_sum[235][11:8] > 6 ? 4'd6 : weighted_sum[235][11:8]);
assign relu_out[236] = (weighted_sum[236][12]==1) ? 4'd0 : (weighted_sum[236][11:8] > 6 ? 4'd6 : weighted_sum[236][11:8]);
assign relu_out[237] = (weighted_sum[237][12]==1) ? 4'd0 : (weighted_sum[237][11:8] > 6 ? 4'd6 : weighted_sum[237][11:8]);
assign relu_out[238] = (weighted_sum[238][12]==1) ? 4'd0 : (weighted_sum[238][11:8] > 6 ? 4'd6 : weighted_sum[238][11:8]);
assign relu_out[239] = (weighted_sum[239][12]==1) ? 4'd0 : (weighted_sum[239][11:8] > 6 ? 4'd6 : weighted_sum[239][11:8]);
assign relu_out[240] = (weighted_sum[240][12]==1) ? 4'd0 : (weighted_sum[240][11:8] > 6 ? 4'd6 : weighted_sum[240][11:8]);
assign relu_out[241] = (weighted_sum[241][12]==1) ? 4'd0 : (weighted_sum[241][11:8] > 6 ? 4'd6 : weighted_sum[241][11:8]);
assign relu_out[242] = (weighted_sum[242][12]==1) ? 4'd0 : (weighted_sum[242][11:8] > 6 ? 4'd6 : weighted_sum[242][11:8]);
assign relu_out[243] = (weighted_sum[243][12]==1) ? 4'd0 : (weighted_sum[243][11:8] > 6 ? 4'd6 : weighted_sum[243][11:8]);
assign relu_out[244] = (weighted_sum[244][12]==1) ? 4'd0 : (weighted_sum[244][11:8] > 6 ? 4'd6 : weighted_sum[244][11:8]);
assign relu_out[245] = (weighted_sum[245][12]==1) ? 4'd0 : (weighted_sum[245][11:8] > 6 ? 4'd6 : weighted_sum[245][11:8]);
assign relu_out[246] = (weighted_sum[246][12]==1) ? 4'd0 : (weighted_sum[246][11:8] > 6 ? 4'd6 : weighted_sum[246][11:8]);
assign relu_out[247] = (weighted_sum[247][12]==1) ? 4'd0 : (weighted_sum[247][11:8] > 6 ? 4'd6 : weighted_sum[247][11:8]);
assign relu_out[248] = (weighted_sum[248][12]==1) ? 4'd0 : (weighted_sum[248][11:8] > 6 ? 4'd6 : weighted_sum[248][11:8]);
assign relu_out[249] = (weighted_sum[249][12]==1) ? 4'd0 : (weighted_sum[249][11:8] > 6 ? 4'd6 : weighted_sum[249][11:8]);
assign relu_out[250] = (weighted_sum[250][12]==1) ? 4'd0 : (weighted_sum[250][11:8] > 6 ? 4'd6 : weighted_sum[250][11:8]);
assign relu_out[251] = (weighted_sum[251][12]==1) ? 4'd0 : (weighted_sum[251][11:8] > 6 ? 4'd6 : weighted_sum[251][11:8]);
assign relu_out[252] = (weighted_sum[252][12]==1) ? 4'd0 : (weighted_sum[252][11:8] > 6 ? 4'd6 : weighted_sum[252][11:8]);
assign relu_out[253] = (weighted_sum[253][12]==1) ? 4'd0 : (weighted_sum[253][11:8] > 6 ? 4'd6 : weighted_sum[253][11:8]);
assign relu_out[254] = (weighted_sum[254][12]==1) ? 4'd0 : (weighted_sum[254][11:8] > 6 ? 4'd6 : weighted_sum[254][11:8]);
assign relu_out[255] = (weighted_sum[255][12]==1) ? 4'd0 : (weighted_sum[255][11:8] > 6 ? 4'd6 : weighted_sum[255][11:8]);
assign relu_out[256] = (weighted_sum[256][12]==1) ? 4'd0 : (weighted_sum[256][11:8] > 6 ? 4'd6 : weighted_sum[256][11:8]);
assign relu_out[257] = (weighted_sum[257][12]==1) ? 4'd0 : (weighted_sum[257][11:8] > 6 ? 4'd6 : weighted_sum[257][11:8]);
assign relu_out[258] = (weighted_sum[258][12]==1) ? 4'd0 : (weighted_sum[258][11:8] > 6 ? 4'd6 : weighted_sum[258][11:8]);
assign relu_out[259] = (weighted_sum[259][12]==1) ? 4'd0 : (weighted_sum[259][11:8] > 6 ? 4'd6 : weighted_sum[259][11:8]);
assign relu_out[260] = (weighted_sum[260][12]==1) ? 4'd0 : (weighted_sum[260][11:8] > 6 ? 4'd6 : weighted_sum[260][11:8]);
assign relu_out[261] = (weighted_sum[261][12]==1) ? 4'd0 : (weighted_sum[261][11:8] > 6 ? 4'd6 : weighted_sum[261][11:8]);
assign relu_out[262] = (weighted_sum[262][12]==1) ? 4'd0 : (weighted_sum[262][11:8] > 6 ? 4'd6 : weighted_sum[262][11:8]);
assign relu_out[263] = (weighted_sum[263][12]==1) ? 4'd0 : (weighted_sum[263][11:8] > 6 ? 4'd6 : weighted_sum[263][11:8]);
assign relu_out[264] = (weighted_sum[264][12]==1) ? 4'd0 : (weighted_sum[264][11:8] > 6 ? 4'd6 : weighted_sum[264][11:8]);
assign relu_out[265] = (weighted_sum[265][12]==1) ? 4'd0 : (weighted_sum[265][11:8] > 6 ? 4'd6 : weighted_sum[265][11:8]);
assign relu_out[266] = (weighted_sum[266][12]==1) ? 4'd0 : (weighted_sum[266][11:8] > 6 ? 4'd6 : weighted_sum[266][11:8]);
assign relu_out[267] = (weighted_sum[267][12]==1) ? 4'd0 : (weighted_sum[267][11:8] > 6 ? 4'd6 : weighted_sum[267][11:8]);
assign relu_out[268] = (weighted_sum[268][12]==1) ? 4'd0 : (weighted_sum[268][11:8] > 6 ? 4'd6 : weighted_sum[268][11:8]);
assign relu_out[269] = (weighted_sum[269][12]==1) ? 4'd0 : (weighted_sum[269][11:8] > 6 ? 4'd6 : weighted_sum[269][11:8]);
assign relu_out[270] = (weighted_sum[270][12]==1) ? 4'd0 : (weighted_sum[270][11:8] > 6 ? 4'd6 : weighted_sum[270][11:8]);
assign relu_out[271] = (weighted_sum[271][12]==1) ? 4'd0 : (weighted_sum[271][11:8] > 6 ? 4'd6 : weighted_sum[271][11:8]);
assign relu_out[272] = (weighted_sum[272][12]==1) ? 4'd0 : (weighted_sum[272][11:8] > 6 ? 4'd6 : weighted_sum[272][11:8]);
assign relu_out[273] = (weighted_sum[273][12]==1) ? 4'd0 : (weighted_sum[273][11:8] > 6 ? 4'd6 : weighted_sum[273][11:8]);
assign relu_out[274] = (weighted_sum[274][12]==1) ? 4'd0 : (weighted_sum[274][11:8] > 6 ? 4'd6 : weighted_sum[274][11:8]);
assign relu_out[275] = (weighted_sum[275][12]==1) ? 4'd0 : (weighted_sum[275][11:8] > 6 ? 4'd6 : weighted_sum[275][11:8]);
assign relu_out[276] = (weighted_sum[276][12]==1) ? 4'd0 : (weighted_sum[276][11:8] > 6 ? 4'd6 : weighted_sum[276][11:8]);
assign relu_out[277] = (weighted_sum[277][12]==1) ? 4'd0 : (weighted_sum[277][11:8] > 6 ? 4'd6 : weighted_sum[277][11:8]);
assign relu_out[278] = (weighted_sum[278][12]==1) ? 4'd0 : (weighted_sum[278][11:8] > 6 ? 4'd6 : weighted_sum[278][11:8]);
assign relu_out[279] = (weighted_sum[279][12]==1) ? 4'd0 : (weighted_sum[279][11:8] > 6 ? 4'd6 : weighted_sum[279][11:8]);
assign relu_out[280] = (weighted_sum[280][12]==1) ? 4'd0 : (weighted_sum[280][11:8] > 6 ? 4'd6 : weighted_sum[280][11:8]);
assign relu_out[281] = (weighted_sum[281][12]==1) ? 4'd0 : (weighted_sum[281][11:8] > 6 ? 4'd6 : weighted_sum[281][11:8]);
assign relu_out[282] = (weighted_sum[282][12]==1) ? 4'd0 : (weighted_sum[282][11:8] > 6 ? 4'd6 : weighted_sum[282][11:8]);
assign relu_out[283] = (weighted_sum[283][12]==1) ? 4'd0 : (weighted_sum[283][11:8] > 6 ? 4'd6 : weighted_sum[283][11:8]);
assign relu_out[284] = (weighted_sum[284][12]==1) ? 4'd0 : (weighted_sum[284][11:8] > 6 ? 4'd6 : weighted_sum[284][11:8]);
assign relu_out[285] = (weighted_sum[285][12]==1) ? 4'd0 : (weighted_sum[285][11:8] > 6 ? 4'd6 : weighted_sum[285][11:8]);
assign relu_out[286] = (weighted_sum[286][12]==1) ? 4'd0 : (weighted_sum[286][11:8] > 6 ? 4'd6 : weighted_sum[286][11:8]);
assign relu_out[287] = (weighted_sum[287][12]==1) ? 4'd0 : (weighted_sum[287][11:8] > 6 ? 4'd6 : weighted_sum[287][11:8]);
assign relu_out[288] = (weighted_sum[288][12]==1) ? 4'd0 : (weighted_sum[288][11:8] > 6 ? 4'd6 : weighted_sum[288][11:8]);
assign relu_out[289] = (weighted_sum[289][12]==1) ? 4'd0 : (weighted_sum[289][11:8] > 6 ? 4'd6 : weighted_sum[289][11:8]);
assign relu_out[290] = (weighted_sum[290][12]==1) ? 4'd0 : (weighted_sum[290][11:8] > 6 ? 4'd6 : weighted_sum[290][11:8]);
assign relu_out[291] = (weighted_sum[291][12]==1) ? 4'd0 : (weighted_sum[291][11:8] > 6 ? 4'd6 : weighted_sum[291][11:8]);
assign relu_out[292] = (weighted_sum[292][12]==1) ? 4'd0 : (weighted_sum[292][11:8] > 6 ? 4'd6 : weighted_sum[292][11:8]);
assign relu_out[293] = (weighted_sum[293][12]==1) ? 4'd0 : (weighted_sum[293][11:8] > 6 ? 4'd6 : weighted_sum[293][11:8]);
assign relu_out[294] = (weighted_sum[294][12]==1) ? 4'd0 : (weighted_sum[294][11:8] > 6 ? 4'd6 : weighted_sum[294][11:8]);
assign relu_out[295] = (weighted_sum[295][12]==1) ? 4'd0 : (weighted_sum[295][11:8] > 6 ? 4'd6 : weighted_sum[295][11:8]);
assign relu_out[296] = (weighted_sum[296][12]==1) ? 4'd0 : (weighted_sum[296][11:8] > 6 ? 4'd6 : weighted_sum[296][11:8]);
assign relu_out[297] = (weighted_sum[297][12]==1) ? 4'd0 : (weighted_sum[297][11:8] > 6 ? 4'd6 : weighted_sum[297][11:8]);
assign relu_out[298] = (weighted_sum[298][12]==1) ? 4'd0 : (weighted_sum[298][11:8] > 6 ? 4'd6 : weighted_sum[298][11:8]);
assign relu_out[299] = (weighted_sum[299][12]==1) ? 4'd0 : (weighted_sum[299][11:8] > 6 ? 4'd6 : weighted_sum[299][11:8]);
assign relu_out[300] = (weighted_sum[300][12]==1) ? 4'd0 : (weighted_sum[300][11:8] > 6 ? 4'd6 : weighted_sum[300][11:8]);
assign relu_out[301] = (weighted_sum[301][12]==1) ? 4'd0 : (weighted_sum[301][11:8] > 6 ? 4'd6 : weighted_sum[301][11:8]);
assign relu_out[302] = (weighted_sum[302][12]==1) ? 4'd0 : (weighted_sum[302][11:8] > 6 ? 4'd6 : weighted_sum[302][11:8]);
assign relu_out[303] = (weighted_sum[303][12]==1) ? 4'd0 : (weighted_sum[303][11:8] > 6 ? 4'd6 : weighted_sum[303][11:8]);
assign relu_out[304] = (weighted_sum[304][12]==1) ? 4'd0 : (weighted_sum[304][11:8] > 6 ? 4'd6 : weighted_sum[304][11:8]);
assign relu_out[305] = (weighted_sum[305][12]==1) ? 4'd0 : (weighted_sum[305][11:8] > 6 ? 4'd6 : weighted_sum[305][11:8]);
assign relu_out[306] = (weighted_sum[306][12]==1) ? 4'd0 : (weighted_sum[306][11:8] > 6 ? 4'd6 : weighted_sum[306][11:8]);
assign relu_out[307] = (weighted_sum[307][12]==1) ? 4'd0 : (weighted_sum[307][11:8] > 6 ? 4'd6 : weighted_sum[307][11:8]);
assign relu_out[308] = (weighted_sum[308][12]==1) ? 4'd0 : (weighted_sum[308][11:8] > 6 ? 4'd6 : weighted_sum[308][11:8]);
assign relu_out[309] = (weighted_sum[309][12]==1) ? 4'd0 : (weighted_sum[309][11:8] > 6 ? 4'd6 : weighted_sum[309][11:8]);
assign relu_out[310] = (weighted_sum[310][12]==1) ? 4'd0 : (weighted_sum[310][11:8] > 6 ? 4'd6 : weighted_sum[310][11:8]);
assign relu_out[311] = (weighted_sum[311][12]==1) ? 4'd0 : (weighted_sum[311][11:8] > 6 ? 4'd6 : weighted_sum[311][11:8]);
assign relu_out[312] = (weighted_sum[312][12]==1) ? 4'd0 : (weighted_sum[312][11:8] > 6 ? 4'd6 : weighted_sum[312][11:8]);
assign relu_out[313] = (weighted_sum[313][12]==1) ? 4'd0 : (weighted_sum[313][11:8] > 6 ? 4'd6 : weighted_sum[313][11:8]);
assign relu_out[314] = (weighted_sum[314][12]==1) ? 4'd0 : (weighted_sum[314][11:8] > 6 ? 4'd6 : weighted_sum[314][11:8]);
assign relu_out[315] = (weighted_sum[315][12]==1) ? 4'd0 : (weighted_sum[315][11:8] > 6 ? 4'd6 : weighted_sum[315][11:8]);
assign relu_out[316] = (weighted_sum[316][12]==1) ? 4'd0 : (weighted_sum[316][11:8] > 6 ? 4'd6 : weighted_sum[316][11:8]);
assign relu_out[317] = (weighted_sum[317][12]==1) ? 4'd0 : (weighted_sum[317][11:8] > 6 ? 4'd6 : weighted_sum[317][11:8]);
assign relu_out[318] = (weighted_sum[318][12]==1) ? 4'd0 : (weighted_sum[318][11:8] > 6 ? 4'd6 : weighted_sum[318][11:8]);
assign relu_out[319] = (weighted_sum[319][12]==1) ? 4'd0 : (weighted_sum[319][11:8] > 6 ? 4'd6 : weighted_sum[319][11:8]);
assign relu_out[320] = (weighted_sum[320][12]==1) ? 4'd0 : (weighted_sum[320][11:8] > 6 ? 4'd6 : weighted_sum[320][11:8]);
assign relu_out[321] = (weighted_sum[321][12]==1) ? 4'd0 : (weighted_sum[321][11:8] > 6 ? 4'd6 : weighted_sum[321][11:8]);
assign relu_out[322] = (weighted_sum[322][12]==1) ? 4'd0 : (weighted_sum[322][11:8] > 6 ? 4'd6 : weighted_sum[322][11:8]);
assign relu_out[323] = (weighted_sum[323][12]==1) ? 4'd0 : (weighted_sum[323][11:8] > 6 ? 4'd6 : weighted_sum[323][11:8]);
assign relu_out[324] = (weighted_sum[324][12]==1) ? 4'd0 : (weighted_sum[324][11:8] > 6 ? 4'd6 : weighted_sum[324][11:8]);
assign relu_out[325] = (weighted_sum[325][12]==1) ? 4'd0 : (weighted_sum[325][11:8] > 6 ? 4'd6 : weighted_sum[325][11:8]);
assign relu_out[326] = (weighted_sum[326][12]==1) ? 4'd0 : (weighted_sum[326][11:8] > 6 ? 4'd6 : weighted_sum[326][11:8]);
assign relu_out[327] = (weighted_sum[327][12]==1) ? 4'd0 : (weighted_sum[327][11:8] > 6 ? 4'd6 : weighted_sum[327][11:8]);
assign relu_out[328] = (weighted_sum[328][12]==1) ? 4'd0 : (weighted_sum[328][11:8] > 6 ? 4'd6 : weighted_sum[328][11:8]);
assign relu_out[329] = (weighted_sum[329][12]==1) ? 4'd0 : (weighted_sum[329][11:8] > 6 ? 4'd6 : weighted_sum[329][11:8]);
assign relu_out[330] = (weighted_sum[330][12]==1) ? 4'd0 : (weighted_sum[330][11:8] > 6 ? 4'd6 : weighted_sum[330][11:8]);
assign relu_out[331] = (weighted_sum[331][12]==1) ? 4'd0 : (weighted_sum[331][11:8] > 6 ? 4'd6 : weighted_sum[331][11:8]);
assign relu_out[332] = (weighted_sum[332][12]==1) ? 4'd0 : (weighted_sum[332][11:8] > 6 ? 4'd6 : weighted_sum[332][11:8]);
assign relu_out[333] = (weighted_sum[333][12]==1) ? 4'd0 : (weighted_sum[333][11:8] > 6 ? 4'd6 : weighted_sum[333][11:8]);
assign relu_out[334] = (weighted_sum[334][12]==1) ? 4'd0 : (weighted_sum[334][11:8] > 6 ? 4'd6 : weighted_sum[334][11:8]);
assign relu_out[335] = (weighted_sum[335][12]==1) ? 4'd0 : (weighted_sum[335][11:8] > 6 ? 4'd6 : weighted_sum[335][11:8]);
assign relu_out[336] = (weighted_sum[336][12]==1) ? 4'd0 : (weighted_sum[336][11:8] > 6 ? 4'd6 : weighted_sum[336][11:8]);
assign relu_out[337] = (weighted_sum[337][12]==1) ? 4'd0 : (weighted_sum[337][11:8] > 6 ? 4'd6 : weighted_sum[337][11:8]);
assign relu_out[338] = (weighted_sum[338][12]==1) ? 4'd0 : (weighted_sum[338][11:8] > 6 ? 4'd6 : weighted_sum[338][11:8]);
assign relu_out[339] = (weighted_sum[339][12]==1) ? 4'd0 : (weighted_sum[339][11:8] > 6 ? 4'd6 : weighted_sum[339][11:8]);
assign relu_out[340] = (weighted_sum[340][12]==1) ? 4'd0 : (weighted_sum[340][11:8] > 6 ? 4'd6 : weighted_sum[340][11:8]);
assign relu_out[341] = (weighted_sum[341][12]==1) ? 4'd0 : (weighted_sum[341][11:8] > 6 ? 4'd6 : weighted_sum[341][11:8]);
assign relu_out[342] = (weighted_sum[342][12]==1) ? 4'd0 : (weighted_sum[342][11:8] > 6 ? 4'd6 : weighted_sum[342][11:8]);
assign relu_out[343] = (weighted_sum[343][12]==1) ? 4'd0 : (weighted_sum[343][11:8] > 6 ? 4'd6 : weighted_sum[343][11:8]);
assign relu_out[344] = (weighted_sum[344][12]==1) ? 4'd0 : (weighted_sum[344][11:8] > 6 ? 4'd6 : weighted_sum[344][11:8]);
assign relu_out[345] = (weighted_sum[345][12]==1) ? 4'd0 : (weighted_sum[345][11:8] > 6 ? 4'd6 : weighted_sum[345][11:8]);
assign relu_out[346] = (weighted_sum[346][12]==1) ? 4'd0 : (weighted_sum[346][11:8] > 6 ? 4'd6 : weighted_sum[346][11:8]);
assign relu_out[347] = (weighted_sum[347][12]==1) ? 4'd0 : (weighted_sum[347][11:8] > 6 ? 4'd6 : weighted_sum[347][11:8]);
assign relu_out[348] = (weighted_sum[348][12]==1) ? 4'd0 : (weighted_sum[348][11:8] > 6 ? 4'd6 : weighted_sum[348][11:8]);
assign relu_out[349] = (weighted_sum[349][12]==1) ? 4'd0 : (weighted_sum[349][11:8] > 6 ? 4'd6 : weighted_sum[349][11:8]);
assign relu_out[350] = (weighted_sum[350][12]==1) ? 4'd0 : (weighted_sum[350][11:8] > 6 ? 4'd6 : weighted_sum[350][11:8]);
assign relu_out[351] = (weighted_sum[351][12]==1) ? 4'd0 : (weighted_sum[351][11:8] > 6 ? 4'd6 : weighted_sum[351][11:8]);
assign relu_out[352] = (weighted_sum[352][12]==1) ? 4'd0 : (weighted_sum[352][11:8] > 6 ? 4'd6 : weighted_sum[352][11:8]);
assign relu_out[353] = (weighted_sum[353][12]==1) ? 4'd0 : (weighted_sum[353][11:8] > 6 ? 4'd6 : weighted_sum[353][11:8]);
assign relu_out[354] = (weighted_sum[354][12]==1) ? 4'd0 : (weighted_sum[354][11:8] > 6 ? 4'd6 : weighted_sum[354][11:8]);
assign relu_out[355] = (weighted_sum[355][12]==1) ? 4'd0 : (weighted_sum[355][11:8] > 6 ? 4'd6 : weighted_sum[355][11:8]);
assign relu_out[356] = (weighted_sum[356][12]==1) ? 4'd0 : (weighted_sum[356][11:8] > 6 ? 4'd6 : weighted_sum[356][11:8]);
assign relu_out[357] = (weighted_sum[357][12]==1) ? 4'd0 : (weighted_sum[357][11:8] > 6 ? 4'd6 : weighted_sum[357][11:8]);
assign relu_out[358] = (weighted_sum[358][12]==1) ? 4'd0 : (weighted_sum[358][11:8] > 6 ? 4'd6 : weighted_sum[358][11:8]);
assign relu_out[359] = (weighted_sum[359][12]==1) ? 4'd0 : (weighted_sum[359][11:8] > 6 ? 4'd6 : weighted_sum[359][11:8]);
assign relu_out[360] = (weighted_sum[360][12]==1) ? 4'd0 : (weighted_sum[360][11:8] > 6 ? 4'd6 : weighted_sum[360][11:8]);
assign relu_out[361] = (weighted_sum[361][12]==1) ? 4'd0 : (weighted_sum[361][11:8] > 6 ? 4'd6 : weighted_sum[361][11:8]);
assign relu_out[362] = (weighted_sum[362][12]==1) ? 4'd0 : (weighted_sum[362][11:8] > 6 ? 4'd6 : weighted_sum[362][11:8]);
assign relu_out[363] = (weighted_sum[363][12]==1) ? 4'd0 : (weighted_sum[363][11:8] > 6 ? 4'd6 : weighted_sum[363][11:8]);
assign relu_out[364] = (weighted_sum[364][12]==1) ? 4'd0 : (weighted_sum[364][11:8] > 6 ? 4'd6 : weighted_sum[364][11:8]);
assign relu_out[365] = (weighted_sum[365][12]==1) ? 4'd0 : (weighted_sum[365][11:8] > 6 ? 4'd6 : weighted_sum[365][11:8]);
assign relu_out[366] = (weighted_sum[366][12]==1) ? 4'd0 : (weighted_sum[366][11:8] > 6 ? 4'd6 : weighted_sum[366][11:8]);
assign relu_out[367] = (weighted_sum[367][12]==1) ? 4'd0 : (weighted_sum[367][11:8] > 6 ? 4'd6 : weighted_sum[367][11:8]);
assign relu_out[368] = (weighted_sum[368][12]==1) ? 4'd0 : (weighted_sum[368][11:8] > 6 ? 4'd6 : weighted_sum[368][11:8]);
assign relu_out[369] = (weighted_sum[369][12]==1) ? 4'd0 : (weighted_sum[369][11:8] > 6 ? 4'd6 : weighted_sum[369][11:8]);
assign relu_out[370] = (weighted_sum[370][12]==1) ? 4'd0 : (weighted_sum[370][11:8] > 6 ? 4'd6 : weighted_sum[370][11:8]);
assign relu_out[371] = (weighted_sum[371][12]==1) ? 4'd0 : (weighted_sum[371][11:8] > 6 ? 4'd6 : weighted_sum[371][11:8]);
assign relu_out[372] = (weighted_sum[372][12]==1) ? 4'd0 : (weighted_sum[372][11:8] > 6 ? 4'd6 : weighted_sum[372][11:8]);
assign relu_out[373] = (weighted_sum[373][12]==1) ? 4'd0 : (weighted_sum[373][11:8] > 6 ? 4'd6 : weighted_sum[373][11:8]);
assign relu_out[374] = (weighted_sum[374][12]==1) ? 4'd0 : (weighted_sum[374][11:8] > 6 ? 4'd6 : weighted_sum[374][11:8]);
assign relu_out[375] = (weighted_sum[375][12]==1) ? 4'd0 : (weighted_sum[375][11:8] > 6 ? 4'd6 : weighted_sum[375][11:8]);
assign relu_out[376] = (weighted_sum[376][12]==1) ? 4'd0 : (weighted_sum[376][11:8] > 6 ? 4'd6 : weighted_sum[376][11:8]);
assign relu_out[377] = (weighted_sum[377][12]==1) ? 4'd0 : (weighted_sum[377][11:8] > 6 ? 4'd6 : weighted_sum[377][11:8]);
assign relu_out[378] = (weighted_sum[378][12]==1) ? 4'd0 : (weighted_sum[378][11:8] > 6 ? 4'd6 : weighted_sum[378][11:8]);
assign relu_out[379] = (weighted_sum[379][12]==1) ? 4'd0 : (weighted_sum[379][11:8] > 6 ? 4'd6 : weighted_sum[379][11:8]);
assign relu_out[380] = (weighted_sum[380][12]==1) ? 4'd0 : (weighted_sum[380][11:8] > 6 ? 4'd6 : weighted_sum[380][11:8]);
assign relu_out[381] = (weighted_sum[381][12]==1) ? 4'd0 : (weighted_sum[381][11:8] > 6 ? 4'd6 : weighted_sum[381][11:8]);
assign relu_out[382] = (weighted_sum[382][12]==1) ? 4'd0 : (weighted_sum[382][11:8] > 6 ? 4'd6 : weighted_sum[382][11:8]);
assign relu_out[383] = (weighted_sum[383][12]==1) ? 4'd0 : (weighted_sum[383][11:8] > 6 ? 4'd6 : weighted_sum[383][11:8]);
assign relu_out[384] = (weighted_sum[384][12]==1) ? 4'd0 : (weighted_sum[384][11:8] > 6 ? 4'd6 : weighted_sum[384][11:8]);
assign relu_out[385] = (weighted_sum[385][12]==1) ? 4'd0 : (weighted_sum[385][11:8] > 6 ? 4'd6 : weighted_sum[385][11:8]);
assign relu_out[386] = (weighted_sum[386][12]==1) ? 4'd0 : (weighted_sum[386][11:8] > 6 ? 4'd6 : weighted_sum[386][11:8]);
assign relu_out[387] = (weighted_sum[387][12]==1) ? 4'd0 : (weighted_sum[387][11:8] > 6 ? 4'd6 : weighted_sum[387][11:8]);
assign relu_out[388] = (weighted_sum[388][12]==1) ? 4'd0 : (weighted_sum[388][11:8] > 6 ? 4'd6 : weighted_sum[388][11:8]);
assign relu_out[389] = (weighted_sum[389][12]==1) ? 4'd0 : (weighted_sum[389][11:8] > 6 ? 4'd6 : weighted_sum[389][11:8]);
assign relu_out[390] = (weighted_sum[390][12]==1) ? 4'd0 : (weighted_sum[390][11:8] > 6 ? 4'd6 : weighted_sum[390][11:8]);
assign relu_out[391] = (weighted_sum[391][12]==1) ? 4'd0 : (weighted_sum[391][11:8] > 6 ? 4'd6 : weighted_sum[391][11:8]);
assign relu_out[392] = (weighted_sum[392][12]==1) ? 4'd0 : (weighted_sum[392][11:8] > 6 ? 4'd6 : weighted_sum[392][11:8]);
assign relu_out[393] = (weighted_sum[393][12]==1) ? 4'd0 : (weighted_sum[393][11:8] > 6 ? 4'd6 : weighted_sum[393][11:8]);
assign relu_out[394] = (weighted_sum[394][12]==1) ? 4'd0 : (weighted_sum[394][11:8] > 6 ? 4'd6 : weighted_sum[394][11:8]);
assign relu_out[395] = (weighted_sum[395][12]==1) ? 4'd0 : (weighted_sum[395][11:8] > 6 ? 4'd6 : weighted_sum[395][11:8]);
assign relu_out[396] = (weighted_sum[396][12]==1) ? 4'd0 : (weighted_sum[396][11:8] > 6 ? 4'd6 : weighted_sum[396][11:8]);
assign relu_out[397] = (weighted_sum[397][12]==1) ? 4'd0 : (weighted_sum[397][11:8] > 6 ? 4'd6 : weighted_sum[397][11:8]);
assign relu_out[398] = (weighted_sum[398][12]==1) ? 4'd0 : (weighted_sum[398][11:8] > 6 ? 4'd6 : weighted_sum[398][11:8]);
assign relu_out[399] = (weighted_sum[399][12]==1) ? 4'd0 : (weighted_sum[399][11:8] > 6 ? 4'd6 : weighted_sum[399][11:8]);
assign relu_out[400] = (weighted_sum[400][12]==1) ? 4'd0 : (weighted_sum[400][11:8] > 6 ? 4'd6 : weighted_sum[400][11:8]);
assign relu_out[401] = (weighted_sum[401][12]==1) ? 4'd0 : (weighted_sum[401][11:8] > 6 ? 4'd6 : weighted_sum[401][11:8]);
assign relu_out[402] = (weighted_sum[402][12]==1) ? 4'd0 : (weighted_sum[402][11:8] > 6 ? 4'd6 : weighted_sum[402][11:8]);
assign relu_out[403] = (weighted_sum[403][12]==1) ? 4'd0 : (weighted_sum[403][11:8] > 6 ? 4'd6 : weighted_sum[403][11:8]);
assign relu_out[404] = (weighted_sum[404][12]==1) ? 4'd0 : (weighted_sum[404][11:8] > 6 ? 4'd6 : weighted_sum[404][11:8]);
assign relu_out[405] = (weighted_sum[405][12]==1) ? 4'd0 : (weighted_sum[405][11:8] > 6 ? 4'd6 : weighted_sum[405][11:8]);
assign relu_out[406] = (weighted_sum[406][12]==1) ? 4'd0 : (weighted_sum[406][11:8] > 6 ? 4'd6 : weighted_sum[406][11:8]);
assign relu_out[407] = (weighted_sum[407][12]==1) ? 4'd0 : (weighted_sum[407][11:8] > 6 ? 4'd6 : weighted_sum[407][11:8]);
assign relu_out[408] = (weighted_sum[408][12]==1) ? 4'd0 : (weighted_sum[408][11:8] > 6 ? 4'd6 : weighted_sum[408][11:8]);
assign relu_out[409] = (weighted_sum[409][12]==1) ? 4'd0 : (weighted_sum[409][11:8] > 6 ? 4'd6 : weighted_sum[409][11:8]);
assign relu_out[410] = (weighted_sum[410][12]==1) ? 4'd0 : (weighted_sum[410][11:8] > 6 ? 4'd6 : weighted_sum[410][11:8]);
assign relu_out[411] = (weighted_sum[411][12]==1) ? 4'd0 : (weighted_sum[411][11:8] > 6 ? 4'd6 : weighted_sum[411][11:8]);
assign relu_out[412] = (weighted_sum[412][12]==1) ? 4'd0 : (weighted_sum[412][11:8] > 6 ? 4'd6 : weighted_sum[412][11:8]);
assign relu_out[413] = (weighted_sum[413][12]==1) ? 4'd0 : (weighted_sum[413][11:8] > 6 ? 4'd6 : weighted_sum[413][11:8]);
assign relu_out[414] = (weighted_sum[414][12]==1) ? 4'd0 : (weighted_sum[414][11:8] > 6 ? 4'd6 : weighted_sum[414][11:8]);
assign relu_out[415] = (weighted_sum[415][12]==1) ? 4'd0 : (weighted_sum[415][11:8] > 6 ? 4'd6 : weighted_sum[415][11:8]);
assign relu_out[416] = (weighted_sum[416][12]==1) ? 4'd0 : (weighted_sum[416][11:8] > 6 ? 4'd6 : weighted_sum[416][11:8]);
assign relu_out[417] = (weighted_sum[417][12]==1) ? 4'd0 : (weighted_sum[417][11:8] > 6 ? 4'd6 : weighted_sum[417][11:8]);
assign relu_out[418] = (weighted_sum[418][12]==1) ? 4'd0 : (weighted_sum[418][11:8] > 6 ? 4'd6 : weighted_sum[418][11:8]);
assign relu_out[419] = (weighted_sum[419][12]==1) ? 4'd0 : (weighted_sum[419][11:8] > 6 ? 4'd6 : weighted_sum[419][11:8]);
assign relu_out[420] = (weighted_sum[420][12]==1) ? 4'd0 : (weighted_sum[420][11:8] > 6 ? 4'd6 : weighted_sum[420][11:8]);
assign relu_out[421] = (weighted_sum[421][12]==1) ? 4'd0 : (weighted_sum[421][11:8] > 6 ? 4'd6 : weighted_sum[421][11:8]);
assign relu_out[422] = (weighted_sum[422][12]==1) ? 4'd0 : (weighted_sum[422][11:8] > 6 ? 4'd6 : weighted_sum[422][11:8]);
assign relu_out[423] = (weighted_sum[423][12]==1) ? 4'd0 : (weighted_sum[423][11:8] > 6 ? 4'd6 : weighted_sum[423][11:8]);
assign relu_out[424] = (weighted_sum[424][12]==1) ? 4'd0 : (weighted_sum[424][11:8] > 6 ? 4'd6 : weighted_sum[424][11:8]);
assign relu_out[425] = (weighted_sum[425][12]==1) ? 4'd0 : (weighted_sum[425][11:8] > 6 ? 4'd6 : weighted_sum[425][11:8]);
assign relu_out[426] = (weighted_sum[426][12]==1) ? 4'd0 : (weighted_sum[426][11:8] > 6 ? 4'd6 : weighted_sum[426][11:8]);
assign relu_out[427] = (weighted_sum[427][12]==1) ? 4'd0 : (weighted_sum[427][11:8] > 6 ? 4'd6 : weighted_sum[427][11:8]);
assign relu_out[428] = (weighted_sum[428][12]==1) ? 4'd0 : (weighted_sum[428][11:8] > 6 ? 4'd6 : weighted_sum[428][11:8]);
assign relu_out[429] = (weighted_sum[429][12]==1) ? 4'd0 : (weighted_sum[429][11:8] > 6 ? 4'd6 : weighted_sum[429][11:8]);
assign relu_out[430] = (weighted_sum[430][12]==1) ? 4'd0 : (weighted_sum[430][11:8] > 6 ? 4'd6 : weighted_sum[430][11:8]);
assign relu_out[431] = (weighted_sum[431][12]==1) ? 4'd0 : (weighted_sum[431][11:8] > 6 ? 4'd6 : weighted_sum[431][11:8]);
assign relu_out[432] = (weighted_sum[432][12]==1) ? 4'd0 : (weighted_sum[432][11:8] > 6 ? 4'd6 : weighted_sum[432][11:8]);
assign relu_out[433] = (weighted_sum[433][12]==1) ? 4'd0 : (weighted_sum[433][11:8] > 6 ? 4'd6 : weighted_sum[433][11:8]);
assign relu_out[434] = (weighted_sum[434][12]==1) ? 4'd0 : (weighted_sum[434][11:8] > 6 ? 4'd6 : weighted_sum[434][11:8]);
assign relu_out[435] = (weighted_sum[435][12]==1) ? 4'd0 : (weighted_sum[435][11:8] > 6 ? 4'd6 : weighted_sum[435][11:8]);
assign relu_out[436] = (weighted_sum[436][12]==1) ? 4'd0 : (weighted_sum[436][11:8] > 6 ? 4'd6 : weighted_sum[436][11:8]);
assign relu_out[437] = (weighted_sum[437][12]==1) ? 4'd0 : (weighted_sum[437][11:8] > 6 ? 4'd6 : weighted_sum[437][11:8]);
assign relu_out[438] = (weighted_sum[438][12]==1) ? 4'd0 : (weighted_sum[438][11:8] > 6 ? 4'd6 : weighted_sum[438][11:8]);
assign relu_out[439] = (weighted_sum[439][12]==1) ? 4'd0 : (weighted_sum[439][11:8] > 6 ? 4'd6 : weighted_sum[439][11:8]);
assign relu_out[440] = (weighted_sum[440][12]==1) ? 4'd0 : (weighted_sum[440][11:8] > 6 ? 4'd6 : weighted_sum[440][11:8]);
assign relu_out[441] = (weighted_sum[441][12]==1) ? 4'd0 : (weighted_sum[441][11:8] > 6 ? 4'd6 : weighted_sum[441][11:8]);
assign relu_out[442] = (weighted_sum[442][12]==1) ? 4'd0 : (weighted_sum[442][11:8] > 6 ? 4'd6 : weighted_sum[442][11:8]);
assign relu_out[443] = (weighted_sum[443][12]==1) ? 4'd0 : (weighted_sum[443][11:8] > 6 ? 4'd6 : weighted_sum[443][11:8]);
assign relu_out[444] = (weighted_sum[444][12]==1) ? 4'd0 : (weighted_sum[444][11:8] > 6 ? 4'd6 : weighted_sum[444][11:8]);
assign relu_out[445] = (weighted_sum[445][12]==1) ? 4'd0 : (weighted_sum[445][11:8] > 6 ? 4'd6 : weighted_sum[445][11:8]);
assign relu_out[446] = (weighted_sum[446][12]==1) ? 4'd0 : (weighted_sum[446][11:8] > 6 ? 4'd6 : weighted_sum[446][11:8]);
assign relu_out[447] = (weighted_sum[447][12]==1) ? 4'd0 : (weighted_sum[447][11:8] > 6 ? 4'd6 : weighted_sum[447][11:8]);
assign relu_out[448] = (weighted_sum[448][12]==1) ? 4'd0 : (weighted_sum[448][11:8] > 6 ? 4'd6 : weighted_sum[448][11:8]);
assign relu_out[449] = (weighted_sum[449][12]==1) ? 4'd0 : (weighted_sum[449][11:8] > 6 ? 4'd6 : weighted_sum[449][11:8]);
assign relu_out[450] = (weighted_sum[450][12]==1) ? 4'd0 : (weighted_sum[450][11:8] > 6 ? 4'd6 : weighted_sum[450][11:8]);
assign relu_out[451] = (weighted_sum[451][12]==1) ? 4'd0 : (weighted_sum[451][11:8] > 6 ? 4'd6 : weighted_sum[451][11:8]);
assign relu_out[452] = (weighted_sum[452][12]==1) ? 4'd0 : (weighted_sum[452][11:8] > 6 ? 4'd6 : weighted_sum[452][11:8]);
assign relu_out[453] = (weighted_sum[453][12]==1) ? 4'd0 : (weighted_sum[453][11:8] > 6 ? 4'd6 : weighted_sum[453][11:8]);
assign relu_out[454] = (weighted_sum[454][12]==1) ? 4'd0 : (weighted_sum[454][11:8] > 6 ? 4'd6 : weighted_sum[454][11:8]);
assign relu_out[455] = (weighted_sum[455][12]==1) ? 4'd0 : (weighted_sum[455][11:8] > 6 ? 4'd6 : weighted_sum[455][11:8]);
assign relu_out[456] = (weighted_sum[456][12]==1) ? 4'd0 : (weighted_sum[456][11:8] > 6 ? 4'd6 : weighted_sum[456][11:8]);
assign relu_out[457] = (weighted_sum[457][12]==1) ? 4'd0 : (weighted_sum[457][11:8] > 6 ? 4'd6 : weighted_sum[457][11:8]);
assign relu_out[458] = (weighted_sum[458][12]==1) ? 4'd0 : (weighted_sum[458][11:8] > 6 ? 4'd6 : weighted_sum[458][11:8]);
assign relu_out[459] = (weighted_sum[459][12]==1) ? 4'd0 : (weighted_sum[459][11:8] > 6 ? 4'd6 : weighted_sum[459][11:8]);
assign relu_out[460] = (weighted_sum[460][12]==1) ? 4'd0 : (weighted_sum[460][11:8] > 6 ? 4'd6 : weighted_sum[460][11:8]);
assign relu_out[461] = (weighted_sum[461][12]==1) ? 4'd0 : (weighted_sum[461][11:8] > 6 ? 4'd6 : weighted_sum[461][11:8]);
assign relu_out[462] = (weighted_sum[462][12]==1) ? 4'd0 : (weighted_sum[462][11:8] > 6 ? 4'd6 : weighted_sum[462][11:8]);
assign relu_out[463] = (weighted_sum[463][12]==1) ? 4'd0 : (weighted_sum[463][11:8] > 6 ? 4'd6 : weighted_sum[463][11:8]);
assign relu_out[464] = (weighted_sum[464][12]==1) ? 4'd0 : (weighted_sum[464][11:8] > 6 ? 4'd6 : weighted_sum[464][11:8]);
assign relu_out[465] = (weighted_sum[465][12]==1) ? 4'd0 : (weighted_sum[465][11:8] > 6 ? 4'd6 : weighted_sum[465][11:8]);
assign relu_out[466] = (weighted_sum[466][12]==1) ? 4'd0 : (weighted_sum[466][11:8] > 6 ? 4'd6 : weighted_sum[466][11:8]);
assign relu_out[467] = (weighted_sum[467][12]==1) ? 4'd0 : (weighted_sum[467][11:8] > 6 ? 4'd6 : weighted_sum[467][11:8]);
assign relu_out[468] = (weighted_sum[468][12]==1) ? 4'd0 : (weighted_sum[468][11:8] > 6 ? 4'd6 : weighted_sum[468][11:8]);
assign relu_out[469] = (weighted_sum[469][12]==1) ? 4'd0 : (weighted_sum[469][11:8] > 6 ? 4'd6 : weighted_sum[469][11:8]);
assign relu_out[470] = (weighted_sum[470][12]==1) ? 4'd0 : (weighted_sum[470][11:8] > 6 ? 4'd6 : weighted_sum[470][11:8]);
assign relu_out[471] = (weighted_sum[471][12]==1) ? 4'd0 : (weighted_sum[471][11:8] > 6 ? 4'd6 : weighted_sum[471][11:8]);
assign relu_out[472] = (weighted_sum[472][12]==1) ? 4'd0 : (weighted_sum[472][11:8] > 6 ? 4'd6 : weighted_sum[472][11:8]);
assign relu_out[473] = (weighted_sum[473][12]==1) ? 4'd0 : (weighted_sum[473][11:8] > 6 ? 4'd6 : weighted_sum[473][11:8]);
assign relu_out[474] = (weighted_sum[474][12]==1) ? 4'd0 : (weighted_sum[474][11:8] > 6 ? 4'd6 : weighted_sum[474][11:8]);
assign relu_out[475] = (weighted_sum[475][12]==1) ? 4'd0 : (weighted_sum[475][11:8] > 6 ? 4'd6 : weighted_sum[475][11:8]);
assign relu_out[476] = (weighted_sum[476][12]==1) ? 4'd0 : (weighted_sum[476][11:8] > 6 ? 4'd6 : weighted_sum[476][11:8]);
assign relu_out[477] = (weighted_sum[477][12]==1) ? 4'd0 : (weighted_sum[477][11:8] > 6 ? 4'd6 : weighted_sum[477][11:8]);
assign relu_out[478] = (weighted_sum[478][12]==1) ? 4'd0 : (weighted_sum[478][11:8] > 6 ? 4'd6 : weighted_sum[478][11:8]);
assign relu_out[479] = (weighted_sum[479][12]==1) ? 4'd0 : (weighted_sum[479][11:8] > 6 ? 4'd6 : weighted_sum[479][11:8]);
assign relu_out[480] = (weighted_sum[480][12]==1) ? 4'd0 : (weighted_sum[480][11:8] > 6 ? 4'd6 : weighted_sum[480][11:8]);
assign relu_out[481] = (weighted_sum[481][12]==1) ? 4'd0 : (weighted_sum[481][11:8] > 6 ? 4'd6 : weighted_sum[481][11:8]);
assign relu_out[482] = (weighted_sum[482][12]==1) ? 4'd0 : (weighted_sum[482][11:8] > 6 ? 4'd6 : weighted_sum[482][11:8]);
assign relu_out[483] = (weighted_sum[483][12]==1) ? 4'd0 : (weighted_sum[483][11:8] > 6 ? 4'd6 : weighted_sum[483][11:8]);
assign relu_out[484] = (weighted_sum[484][12]==1) ? 4'd0 : (weighted_sum[484][11:8] > 6 ? 4'd6 : weighted_sum[484][11:8]);
assign relu_out[485] = (weighted_sum[485][12]==1) ? 4'd0 : (weighted_sum[485][11:8] > 6 ? 4'd6 : weighted_sum[485][11:8]);
assign relu_out[486] = (weighted_sum[486][12]==1) ? 4'd0 : (weighted_sum[486][11:8] > 6 ? 4'd6 : weighted_sum[486][11:8]);
assign relu_out[487] = (weighted_sum[487][12]==1) ? 4'd0 : (weighted_sum[487][11:8] > 6 ? 4'd6 : weighted_sum[487][11:8]);
assign relu_out[488] = (weighted_sum[488][12]==1) ? 4'd0 : (weighted_sum[488][11:8] > 6 ? 4'd6 : weighted_sum[488][11:8]);
assign relu_out[489] = (weighted_sum[489][12]==1) ? 4'd0 : (weighted_sum[489][11:8] > 6 ? 4'd6 : weighted_sum[489][11:8]);
assign relu_out[490] = (weighted_sum[490][12]==1) ? 4'd0 : (weighted_sum[490][11:8] > 6 ? 4'd6 : weighted_sum[490][11:8]);
assign relu_out[491] = (weighted_sum[491][12]==1) ? 4'd0 : (weighted_sum[491][11:8] > 6 ? 4'd6 : weighted_sum[491][11:8]);
assign relu_out[492] = (weighted_sum[492][12]==1) ? 4'd0 : (weighted_sum[492][11:8] > 6 ? 4'd6 : weighted_sum[492][11:8]);
assign relu_out[493] = (weighted_sum[493][12]==1) ? 4'd0 : (weighted_sum[493][11:8] > 6 ? 4'd6 : weighted_sum[493][11:8]);
assign relu_out[494] = (weighted_sum[494][12]==1) ? 4'd0 : (weighted_sum[494][11:8] > 6 ? 4'd6 : weighted_sum[494][11:8]);
assign relu_out[495] = (weighted_sum[495][12]==1) ? 4'd0 : (weighted_sum[495][11:8] > 6 ? 4'd6 : weighted_sum[495][11:8]);
assign relu_out[496] = (weighted_sum[496][12]==1) ? 4'd0 : (weighted_sum[496][11:8] > 6 ? 4'd6 : weighted_sum[496][11:8]);
assign relu_out[497] = (weighted_sum[497][12]==1) ? 4'd0 : (weighted_sum[497][11:8] > 6 ? 4'd6 : weighted_sum[497][11:8]);
assign relu_out[498] = (weighted_sum[498][12]==1) ? 4'd0 : (weighted_sum[498][11:8] > 6 ? 4'd6 : weighted_sum[498][11:8]);
assign relu_out[499] = (weighted_sum[499][12]==1) ? 4'd0 : (weighted_sum[499][11:8] > 6 ? 4'd6 : weighted_sum[499][11:8]);
assign relu_out[500] = (weighted_sum[500][12]==1) ? 4'd0 : (weighted_sum[500][11:8] > 6 ? 4'd6 : weighted_sum[500][11:8]);
assign relu_out[501] = (weighted_sum[501][12]==1) ? 4'd0 : (weighted_sum[501][11:8] > 6 ? 4'd6 : weighted_sum[501][11:8]);
assign relu_out[502] = (weighted_sum[502][12]==1) ? 4'd0 : (weighted_sum[502][11:8] > 6 ? 4'd6 : weighted_sum[502][11:8]);
assign relu_out[503] = (weighted_sum[503][12]==1) ? 4'd0 : (weighted_sum[503][11:8] > 6 ? 4'd6 : weighted_sum[503][11:8]);
assign relu_out[504] = (weighted_sum[504][12]==1) ? 4'd0 : (weighted_sum[504][11:8] > 6 ? 4'd6 : weighted_sum[504][11:8]);
assign relu_out[505] = (weighted_sum[505][12]==1) ? 4'd0 : (weighted_sum[505][11:8] > 6 ? 4'd6 : weighted_sum[505][11:8]);
assign relu_out[506] = (weighted_sum[506][12]==1) ? 4'd0 : (weighted_sum[506][11:8] > 6 ? 4'd6 : weighted_sum[506][11:8]);
assign out = {relu_out[506],relu_out[505],relu_out[504],relu_out[503],relu_out[502],relu_out[501],relu_out[500],relu_out[499],relu_out[498],relu_out[497],relu_out[496],relu_out[495],relu_out[494],relu_out[493],relu_out[492],relu_out[491],relu_out[490],relu_out[489],relu_out[488],relu_out[487],relu_out[486],relu_out[485],relu_out[484],relu_out[483],relu_out[482],relu_out[481],relu_out[480],relu_out[479],relu_out[478],relu_out[477],relu_out[476],relu_out[475],relu_out[474],relu_out[473],relu_out[472],relu_out[471],relu_out[470],relu_out[469],relu_out[468],relu_out[467],relu_out[466],relu_out[465],relu_out[464],relu_out[463],relu_out[462],relu_out[461],relu_out[460],relu_out[459],relu_out[458],relu_out[457],relu_out[456],relu_out[455],relu_out[454],relu_out[453],relu_out[452],relu_out[451],relu_out[450],relu_out[449],relu_out[448],relu_out[447],relu_out[446],relu_out[445],relu_out[444],relu_out[443],relu_out[442],relu_out[441],relu_out[440],relu_out[439],relu_out[438],relu_out[437],relu_out[436],relu_out[435],relu_out[434],relu_out[433],relu_out[432],relu_out[431],relu_out[430],relu_out[429],relu_out[428],relu_out[427],relu_out[426],relu_out[425],relu_out[424],relu_out[423],relu_out[422],relu_out[421],relu_out[420],relu_out[419],relu_out[418],relu_out[417],relu_out[416],relu_out[415],relu_out[414],relu_out[413],relu_out[412],relu_out[411],relu_out[410],relu_out[409],relu_out[408],relu_out[407],relu_out[406],relu_out[405],relu_out[404],relu_out[403],relu_out[402],relu_out[401],relu_out[400],relu_out[399],relu_out[398],relu_out[397],relu_out[396],relu_out[395],relu_out[394],relu_out[393],relu_out[392],relu_out[391],relu_out[390],relu_out[389],relu_out[388],relu_out[387],relu_out[386],relu_out[385],relu_out[384],relu_out[383],relu_out[382],relu_out[381],relu_out[380],relu_out[379],relu_out[378],relu_out[377],relu_out[376],relu_out[375],relu_out[374],relu_out[373],relu_out[372],relu_out[371],relu_out[370],relu_out[369],relu_out[368],relu_out[367],relu_out[366],relu_out[365],relu_out[364],relu_out[363],relu_out[362],relu_out[361],relu_out[360],relu_out[359],relu_out[358],relu_out[357],relu_out[356],relu_out[355],relu_out[354],relu_out[353],relu_out[352],relu_out[351],relu_out[350],relu_out[349],relu_out[348],relu_out[347],relu_out[346],relu_out[345],relu_out[344],relu_out[343],relu_out[342],relu_out[341],relu_out[340],relu_out[339],relu_out[338],relu_out[337],relu_out[336],relu_out[335],relu_out[334],relu_out[333],relu_out[332],relu_out[331],relu_out[330],relu_out[329],relu_out[328],relu_out[327],relu_out[326],relu_out[325],relu_out[324],relu_out[323],relu_out[322],relu_out[321],relu_out[320],relu_out[319],relu_out[318],relu_out[317],relu_out[316],relu_out[315],relu_out[314],relu_out[313],relu_out[312],relu_out[311],relu_out[310],relu_out[309],relu_out[308],relu_out[307],relu_out[306],relu_out[305],relu_out[304],relu_out[303],relu_out[302],relu_out[301],relu_out[300],relu_out[299],relu_out[298],relu_out[297],relu_out[296],relu_out[295],relu_out[294],relu_out[293],relu_out[292],relu_out[291],relu_out[290],relu_out[289],relu_out[288],relu_out[287],relu_out[286],relu_out[285],relu_out[284],relu_out[283],relu_out[282],relu_out[281],relu_out[280],relu_out[279],relu_out[278],relu_out[277],relu_out[276],relu_out[275],relu_out[274],relu_out[273],relu_out[272],relu_out[271],relu_out[270],relu_out[269],relu_out[268],relu_out[267],relu_out[266],relu_out[265],relu_out[264],relu_out[263],relu_out[262],relu_out[261],relu_out[260],relu_out[259],relu_out[258],relu_out[257],relu_out[256],relu_out[255],relu_out[254],relu_out[253],relu_out[252],relu_out[251],relu_out[250],relu_out[249],relu_out[248],relu_out[247],relu_out[246],relu_out[245],relu_out[244],relu_out[243],relu_out[242],relu_out[241],relu_out[240],relu_out[239],relu_out[238],relu_out[237],relu_out[236],relu_out[235],relu_out[234],relu_out[233],relu_out[232],relu_out[231],relu_out[230],relu_out[229],relu_out[228],relu_out[227],relu_out[226],relu_out[225],relu_out[224],relu_out[223],relu_out[222],relu_out[221],relu_out[220],relu_out[219],relu_out[218],relu_out[217],relu_out[216],relu_out[215],relu_out[214],relu_out[213],relu_out[212],relu_out[211],relu_out[210],relu_out[209],relu_out[208],relu_out[207],relu_out[206],relu_out[205],relu_out[204],relu_out[203],relu_out[202],relu_out[201],relu_out[200],relu_out[199],relu_out[198],relu_out[197],relu_out[196],relu_out[195],relu_out[194],relu_out[193],relu_out[192],relu_out[191],relu_out[190],relu_out[189],relu_out[188],relu_out[187],relu_out[186],relu_out[185],relu_out[184],relu_out[183],relu_out[182],relu_out[181],relu_out[180],relu_out[179],relu_out[178],relu_out[177],relu_out[176],relu_out[175],relu_out[174],relu_out[173],relu_out[172],relu_out[171],relu_out[170],relu_out[169],relu_out[168],relu_out[167],relu_out[166],relu_out[165],relu_out[164],relu_out[163],relu_out[162],relu_out[161],relu_out[160],relu_out[159],relu_out[158],relu_out[157],relu_out[156],relu_out[155],relu_out[154],relu_out[153],relu_out[152],relu_out[151],relu_out[150],relu_out[149],relu_out[148],relu_out[147],relu_out[146],relu_out[145],relu_out[144],relu_out[143],relu_out[142],relu_out[141],relu_out[140],relu_out[139],relu_out[138],relu_out[137],relu_out[136],relu_out[135],relu_out[134],relu_out[133],relu_out[132],relu_out[131],relu_out[130],relu_out[129],relu_out[128],relu_out[127],relu_out[126],relu_out[125],relu_out[124],relu_out[123],relu_out[122],relu_out[121],relu_out[120],relu_out[119],relu_out[118],relu_out[117],relu_out[116],relu_out[115],relu_out[114],relu_out[113],relu_out[112],relu_out[111],relu_out[110],relu_out[109],relu_out[108],relu_out[107],relu_out[106],relu_out[105],relu_out[104],relu_out[103],relu_out[102],relu_out[101],relu_out[100],relu_out[99],relu_out[98],relu_out[97],relu_out[96],relu_out[95],relu_out[94],relu_out[93],relu_out[92],relu_out[91],relu_out[90],relu_out[89],relu_out[88],relu_out[87],relu_out[86],relu_out[85],relu_out[84],relu_out[83],relu_out[82],relu_out[81],relu_out[80],relu_out[79],relu_out[78],relu_out[77],relu_out[76],relu_out[75],relu_out[74],relu_out[73],relu_out[72],relu_out[71],relu_out[70],relu_out[69],relu_out[68],relu_out[67],relu_out[66],relu_out[65],relu_out[64],relu_out[63],relu_out[62],relu_out[61],relu_out[60],relu_out[59],relu_out[58],relu_out[57],relu_out[56],relu_out[55],relu_out[54],relu_out[53],relu_out[52],relu_out[51],relu_out[50],relu_out[49],relu_out[48],relu_out[47],relu_out[46],relu_out[45],relu_out[44],relu_out[43],relu_out[42],relu_out[41],relu_out[40],relu_out[39],relu_out[38],relu_out[37],relu_out[36],relu_out[35],relu_out[34],relu_out[33],relu_out[32],relu_out[31],relu_out[30],relu_out[29],relu_out[28],relu_out[27],relu_out[26],relu_out[25],relu_out[24],relu_out[23],relu_out[22],relu_out[21],relu_out[20],relu_out[19],relu_out[18],relu_out[17],relu_out[16],relu_out[15],relu_out[14],relu_out[13],relu_out[12],relu_out[11],relu_out[10],relu_out[9],relu_out[8],relu_out[7],relu_out[6],relu_out[5],relu_out[4],relu_out[3],relu_out[2],relu_out[1],relu_out[0]};

endmodule
