module fc2 (
	input [3:0] in [0:31],
	input clk,
	input rst,
	output [3:0] out [0:31]
);

logic [8:0] weighted_sum [0:31];
logic [8:0] sharing0_r, sharing0_w;
logic [8:0] sharing1_r, sharing1_w;
logic [8:0] sharing2_r, sharing2_w;
logic [8:0] sharing3_r, sharing3_w;
logic [8:0] sharing4_r, sharing4_w;
logic [8:0] sharing5_r, sharing5_w;
logic [8:0] sharing6_r, sharing6_w;
logic [8:0] sharing7_r, sharing7_w;
logic [8:0] sharing8_r, sharing8_w;
logic [8:0] sharing9_r, sharing9_w;
logic [8:0] sharing10_r, sharing10_w;
logic [8:0] sharing11_r, sharing11_w;
logic [8:0] sharing12_r, sharing12_w;
logic [8:0] sharing13_r, sharing13_w;
logic [8:0] sharing14_r, sharing14_w;
logic [8:0] sharing15_r, sharing15_w;
logic [8:0] sharing16_r, sharing16_w;
logic [8:0] sharing17_r, sharing17_w;
logic [8:0] sharing18_r, sharing18_w;
logic [8:0] sharing19_r, sharing19_w;
logic [8:0] sharing20_r, sharing20_w;
logic [8:0] sharing21_r, sharing21_w;
logic [8:0] sharing22_r, sharing22_w;
logic [8:0] sharing23_r, sharing23_w;
logic [8:0] sharing24_r, sharing24_w;
logic [8:0] sharing25_r, sharing25_w;
logic [8:0] sharing26_r, sharing26_w;
logic [8:0] sharing27_r, sharing27_w;
logic [8:0] sharing28_r, sharing28_w;
logic [8:0] sharing29_r, sharing29_w;
logic [8:0] sharing30_r, sharing30_w;
logic [8:0] sharing31_r, sharing31_w;
logic [8:0] sharing32_r, sharing32_w;
logic [8:0] sharing33_r, sharing33_w;
logic [8:0] sharing34_r, sharing34_w;
logic [8:0] sharing35_r, sharing35_w;
logic [8:0] sharing36_r, sharing36_w;
logic [8:0] sharing37_r, sharing37_w;
logic [8:0] sharing38_r, sharing38_w;
logic [8:0] sharing39_r, sharing39_w;
logic [8:0] sharing40_r, sharing40_w;
logic [8:0] sharing41_r, sharing41_w;
logic [8:0] sharing42_r, sharing42_w;
logic [8:0] sharing43_r, sharing43_w;
logic [8:0] sharing44_r, sharing44_w;
logic [8:0] sharing45_r, sharing45_w;
logic [8:0] sharing46_r, sharing46_w;
logic [8:0] sharing47_r, sharing47_w;
logic [8:0] sharing48_r, sharing48_w;
logic [8:0] sharing49_r, sharing49_w;

always_comb begin
	sharing0_w = $signed(in[30])+$signed(-in[26])+$signed(-in[25]);
	sharing1_w = $signed({in[17],1'b0})+$signed({in[7],1'b0})+$signed(-{in[22],1'b0})+$signed(-in[10])+$signed(-in[1])+$signed(-in[31]);
	sharing2_w = $signed(in[25])+$signed(in[2])+$signed({in[3],1'b0})+$signed(in[19])+$signed({in[4],1'b0})+$signed(in[21])+$signed(-{in[21],2'b0})+$signed(-{in[17],1'b0});
	sharing3_w = $signed(in[16])+$signed({in[10],1'b0})+$signed(in[18])+$signed(in[29])+$signed(-{in[26],1'b0})+$signed(-in[11])+$signed(-in[28])+$signed(-in[5])+$signed(-{in[6],2'b0});
	sharing4_w = $signed(in[0])+$signed(in[13])+$signed(-in[8])+$signed(-in[6])+$signed(-in[5])+$signed(-in[29]);
	sharing5_w = $signed({in[18],1'b0})+$signed(in[10])+$signed({in[14],1'b0})+$signed(in[3])+$signed(-{in[23],1'b0})+$signed(-in[11]);
	sharing6_w = $signed(in[18])+$signed(in[26])+$signed(in[3])+$signed(in[23])+$signed(in[7])+$signed(-{in[9],1'b0})+$signed(-{in[26],2'b0})+$signed(-in[28])+$signed(-in[8]);
	sharing7_w = $signed(in[10])+$signed(in[2])+$signed({in[21],1'b0})+$signed(-in[24])+$signed(-{in[17],1'b0})+$signed(-in[25])+$signed(-{in[11],1'b0})+$signed(-{in[14],1'b0})+$signed(-in[6])+$signed(-in[31]);
	sharing8_w = $signed({in[24],1'b0})+$signed({in[10],1'b0})+$signed(in[2])+$signed(in[11])+$signed(in[13])+$signed({in[23],1'b0})+$signed(-in[8])+$signed(-{in[20],1'b0})+$signed(-in[22]);
	sharing9_w = $signed({in[25],1'b0})+$signed(in[9])+$signed(in[1])+$signed(in[3])+$signed(in[28])+$signed(in[7])+$signed(-in[30])+$signed(-in[17]);
	sharing10_w = $signed(in[30])+$signed({in[30],1'b0})+$signed(in[22])+$signed(in[17])+$signed(-in[4])+$signed(-in[15]);
	sharing11_w = $signed({in[19],1'b0})+$signed(in[3])+$signed(-in[1])+$signed(-in[25])+$signed(-{in[18],1'b0})+$signed(-{in[11],1'b0})+$signed(-{in[6],1'b0});
	sharing12_w = $signed(-{in[25],1'b0})+$signed(-in[14])+$signed(-in[26])+$signed(-in[18])+$signed(-in[11])+$signed(-in[3])+$signed(-in[12])+$signed(-in[29])+$signed(-in[5])+$signed(-in[6])+$signed(-in[31]);
	sharing13_w = $signed(in[0])+$signed(in[9])+$signed(in[18])+$signed(in[19])+$signed({in[12],1'b0})+$signed(in[12])+$signed({in[28],1'b0})+$signed({in[6],1'b0})+$signed({in[15],1'b0})+$signed(-in[10])+$signed(-in[20])+$signed(-{in[11],1'b0});
	sharing14_w = $signed(in[14])+$signed(-in[22])+$signed(-in[4])+$signed(-in[31]);
	sharing15_w = $signed(in[28])+$signed(in[12])+$signed({in[13],1'b0})+$signed(in[17])+$signed(-{in[30],1'b0});
	sharing16_w = $signed({in[0],1'b0})+$signed(-{in[24],1'b0})+$signed(-in[9])+$signed(-in[19])+$signed(-{in[31],1'b0})+$signed(-in[15]);
	sharing17_w = $signed({in[0],1'b0})+$signed(in[13])+$signed(in[23])+$signed(in[15])+$signed(-in[16])+$signed(-in[24]);
	sharing18_w = $signed(in[6])+$signed({in[27],1'b0})+$signed(in[7])+$signed(-{in[20],1'b0})+$signed(-{in[25],1'b0})+$signed(-{in[28],1'b0});
	sharing19_w = $signed({in[16],1'b0})+$signed({in[25],1'b0})+$signed(in[2])+$signed({in[20],1'b0})+$signed(in[5])+$signed(in[7])+$signed(-{in[28],1'b0})+$signed(-in[30]);
	sharing20_w = $signed({in[29],1'b0})+$signed(in[13])+$signed(-{in[18],1'b0})+$signed(-in[17])+$signed(-{in[27],1'b0})+$signed(-in[23]);
	sharing21_w = $signed({in[9],1'b0})+$signed(in[17])+$signed(in[25])+$signed(in[3])+$signed({in[20],1'b0})+$signed(in[20])+$signed(-in[8])+$signed(-{in[12],1'b0})+$signed(-in[4])+$signed(-in[31])+$signed(-in[15]);
	sharing22_w = $signed(in[1])+$signed(in[18])+$signed(in[19])+$signed(in[29])+$signed(in[6])+$signed(-in[2]);
	sharing23_w = $signed({in[2],1'b0})+$signed(in[2])+$signed(in[27])+$signed({in[12],1'b0})+$signed(in[22])+$signed(in[31])+$signed(-{in[17],1'b0});
	sharing24_w = $signed({in[3],1'b0})+$signed(in[7])+$signed(-in[0])+$signed(-in[21]);
	sharing25_w = $signed({in[8],1'b0})+$signed(in[16])+$signed(in[24])+$signed(in[26])+$signed(in[27])+$signed({in[28],1'b0})+$signed({in[29],1'b0})+$signed(-{in[2],1'b0})+$signed(-in[14])+$signed(-{in[10],1'b0})+$signed(-{in[31],2'b0});
	sharing26_w = $signed({in[0],1'b0})+$signed(in[30])+$signed(-in[22])+$signed(-in[1]);
	sharing27_w = $signed(in[0])+$signed(in[8])+$signed(in[18])+$signed({in[27],1'b0})+$signed({in[4],2'b0})+$signed(in[12])+$signed({in[23],1'b0})+$signed(in[15])+$signed(-{in[9],1'b0})+$signed(-in[6])+$signed(-{in[25],1'b0})+$signed(-in[13]);
	sharing28_w = $signed({in[5],1'b0})+$signed(-in[10])+$signed(-in[28])+$signed(-in[21])+$signed(-in[31]);
	sharing29_w = $signed({in[10],1'b0})+$signed(in[18])+$signed(in[19])+$signed(in[11])+$signed(in[4])+$signed({in[22],1'b0})+$signed(-in[31])+$signed(-in[23]);
	sharing30_w = $signed(in[0])+$signed(in[24])+$signed(-in[9])+$signed(-{in[12],1'b0})+$signed(-in[28])+$signed(-in[21])+$signed(-in[30])+$signed(-{in[15],1'b0});
	sharing31_w = $signed(in[18])+$signed({in[21],1'b0})+$signed({in[3],1'b0});
	sharing32_w = $signed(in[24])+$signed(-in[20])+$signed(-{in[28],1'b0})+$signed(-in[30])+$signed(-in[1]);
	sharing33_w = $signed({in[5],1'b0})+$signed(in[27])+$signed(-{in[6],3'b0})+$signed(-in[22]);
	sharing34_w = $signed({in[31],1'b0})+$signed(in[9])+$signed(-{in[14],1'b0})+$signed(-{in[21],2'b0});
	sharing35_w = $signed({in[27],1'b0})+$signed({in[14],1'b0})+$signed(in[6])+$signed(in[15])+$signed(in[23])+$signed(-{in[15],2'b0});
	sharing36_w = $signed(in[26])+$signed(in[14])+$signed(-in[0]);
	sharing37_w = $signed(in[11])+$signed(-{in[21],1'b0})+$signed(-in[27]);
	sharing38_w = $signed(in[14])+$signed(in[12])+$signed({in[9],1'b0})+$signed(-{in[11],2'b0});
	sharing39_w = $signed({in[8],1'b0})+$signed(in[20])+$signed(-{in[26],1'b0});
	sharing40_w = $signed(in[12])+$signed(in[27])+$signed(-in[20])+$signed(-in[1]);
	sharing41_w = $signed(in[15])+$signed(-in[19])+$signed(-{in[17],1'b0})+$signed(-in[7]);
	sharing42_w = $signed({in[8],2'b0})+$signed({in[2],1'b0})+$signed(in[28]);
	sharing43_w = $signed({in[24],2'b0})+$signed(-in[14])+$signed(-{in[21],1'b0});
	sharing44_w = $signed({in[17],1'b0})+$signed({in[7],1'b0})+$signed(-{in[27],1'b0})+$signed(-in[5]);
	sharing45_w = $signed({in[16],1'b0})+$signed(in[18])+$signed(-{in[23],1'b0});
	sharing46_w = $signed({in[4],1'b0})+$signed(in[21])+$signed(-{in[9],1'b0});
	sharing47_w = $signed({in[5],2'b0})+$signed({in[21],1'b0})+$signed(-{in[31],2'b0});
	sharing48_w = $signed({in[6],1'b0})+$signed(in[24])+$signed(-{in[5],1'b0});
	sharing49_w = $signed({in[14],1'b0})+$signed({in[26],1'b0})+$signed(in[7]);
end

assign weighted_sum[0] = $signed(-in[24])+$signed(-{in[6],1'b0})+$signed(in[18])+$signed({in[3],1'b0})+$signed(-in[19])+$signed({in[4],2'b0})+$signed(-in[21])+$signed(-{in[14],1'b0})+$signed(-{in[15],3'b0})+$signed({in[15],1'b0})+$signed(sharing0_r)+$signed(sharing1_r)+$signed(sharing42_r)+$signed(1);
assign weighted_sum[1] = $signed(in[8])+$signed({in[1],1'b0})+$signed(-{in[10],2'b0})+$signed(-{in[19],1'b0})+$signed(-{in[12],1'b0})+$signed(in[28])+$signed({in[13],1'b0})+$signed({in[22],1'b0})+$signed(-{in[15],2'b0})+$signed(-in[31])+$signed(sharing17_r)+$signed(-sharing18_r)+$signed(sharing31_r)+$signed(-2);
assign weighted_sum[2] = $signed(-{in[8],2'b0})+$signed(in[8])+$signed(-{in[2],2'b0})+$signed(in[14])+$signed(-{in[12],2'b0})+$signed(-{in[14],3'b0})+$signed({in[22],1'b0})+$signed(-in[30])+$signed(-{in[7],2'b0})+$signed(sharing2_r)+$signed(sharing3_r)+$signed(sharing35_r)+$signed(-4);
assign weighted_sum[3] = $signed({in[0],2'b0})+$signed(-in[16])+$signed({in[25],2'b0})+$signed({in[1],1'b0})+$signed(-in[27])+$signed({in[20],2'b0})+$signed(-in[4])+$signed(-{in[13],2'b0})+$signed(-{in[30],1'b0})+$signed(in[14])+$signed({in[31],2'b0})+$signed({in[15],1'b0})+$signed(sharing4_r)+$signed(sharing5_r)+$signed(0);
assign weighted_sum[4] = $signed({in[0],1'b0})+$signed({in[1],2'b0})+$signed(in[22])+$signed({in[27],1'b0})+$signed(in[19])+$signed(-{in[13],1'b0})+$signed(in[29])+$signed(-in[30])+$signed(in[15])+$signed(sharing6_r)+$signed(sharing7_r)+$signed(-4);
assign weighted_sum[5] = $signed({in[9],1'b0})+$signed(-{in[18],2'b0})+$signed(-{in[27],3'b0})+$signed({in[19],1'b0})+$signed(in[6])+$signed(-in[15])+$signed(-in[23])+$signed(in[31])+$signed(sharing25_r)+$signed(-sharing26_r)+$signed(sharing31_r)+$signed(-sharing44_r)+$signed(2);
assign weighted_sum[6] = $signed({in[2],1'b0})+$signed(-{in[26],1'b0})+$signed(in[28])+$signed(-in[12])+$signed({in[13],1'b0})+$signed({in[22],2'b0})+$signed(in[31])+$signed(sharing4_r)+$signed(-sharing5_r)+$signed(-sharing32_r)+$signed(sharing41_r)+$signed(-sharing46_r)+$signed(-3);
assign weighted_sum[7] = $signed({in[8],1'b0})+$signed({in[24],1'b0})+$signed(in[25])+$signed(-in[6])+$signed({in[12],1'b0})+$signed(-in[4])+$signed({in[7],1'b0})+$signed(-{in[22],2'b0})+$signed(in[22])+$signed(-{in[23],2'b0})+$signed({in[15],1'b0})+$signed(sharing19_r)+$signed(-sharing20_r)+$signed(sharing36_r)+$signed(-sharing37_r)+$signed(1);
assign weighted_sum[8] = $signed(-{in[0],2'b0})+$signed({in[2],1'b0})+$signed(in[18])+$signed({in[27],2'b0})+$signed(-{in[3],2'b0})+$signed({in[12],1'b0})+$signed(-in[4])+$signed({in[28],1'b0})+$signed(in[5])+$signed(-{in[7],2'b0})+$signed({in[31],1'b0})+$signed(sharing8_r)+$signed(sharing9_r)+$signed(sharing43_r)+$signed(2);
assign weighted_sum[9] = $signed({in[24],1'b0})+$signed(in[24])+$signed(in[26])+$signed(in[27])+$signed(-{in[28],1'b0})+$signed({in[5],2'b0})+$signed(-in[21])+$signed(in[29])+$signed({in[14],2'b0})+$signed({in[22],1'b0})+$signed({in[7],2'b0})+$signed(in[23])+$signed(sharing10_r)+$signed(sharing11_r)+$signed(-2);
assign weighted_sum[10] = $signed(in[16])+$signed(in[10])+$signed(-in[27])+$signed(-in[21])+$signed(-in[22])+$signed(sharing12_r)+$signed(sharing32_r)+$signed(-2);
assign weighted_sum[11] = $signed({in[30],1'b0})+$signed(-in[10])+$signed(in[13])+$signed(-in[21])+$signed(sharing21_r)+$signed(-sharing22_r)+$signed(sharing44_r)+$signed(sharing49_r)+$signed(-2);
assign weighted_sum[12] = $signed(-{in[24],1'b0})+$signed(in[8])+$signed(in[6])+$signed(-{in[19],2'b0})+$signed(in[3])+$signed(-{in[5],1'b0})+$signed(-in[13])+$signed(-in[30])+$signed(in[23])+$signed(sharing13_r)+$signed(sharing14_r)+$signed(sharing42_r)+$signed(sharing49_r)+$signed(3);
assign weighted_sum[13] = $signed(in[8])+$signed(-{in[2],2'b0})+$signed(in[26])+$signed(-in[10])+$signed({in[27],1'b0})+$signed(-in[11])+$signed(-{in[12],2'b0})+$signed({in[28],1'b0})+$signed(in[20])+$signed(in[29])+$signed({in[6],1'b0})+$signed(sharing15_r)+$signed(sharing16_r)+$signed(sharing33_r)+$signed(sharing45_r)+$signed(-2);
assign weighted_sum[14] = $signed(-{in[17],2'b0})+$signed({in[25],1'b0})+$signed(in[17])+$signed(-{in[18],2'b0})+$signed(-{in[3],2'b0})+$signed({in[27],1'b0})+$signed(in[3])+$signed(-{in[4],2'b0})+$signed({in[5],1'b0})+$signed(-in[29])+$signed({in[21],1'b0})+$signed({in[6],1'b0})+$signed(-in[14])+$signed(-in[7])+$signed(sharing29_r)+$signed(-sharing30_r)+$signed(0);
assign weighted_sum[15] = $signed(in[0])+$signed({in[1],1'b0})+$signed(-{in[11],3'b0})+$signed({in[20],1'b0})+$signed(-in[4])+$signed(in[5])+$signed(-{in[5],2'b0})+$signed(-in[13])+$signed({in[22],1'b0})+$signed(sharing6_r)+$signed(-sharing7_r)+$signed(-sharing40_r)+$signed(0);
assign weighted_sum[16] = $signed(in[0])+$signed(-{in[1],2'b0})+$signed(in[1])+$signed(-in[26])+$signed(in[11])+$signed(in[19])+$signed(-in[12])+$signed(sharing17_r)+$signed(sharing18_r)+$signed(sharing33_r)+$signed(sharing46_r)+$signed(0);
assign weighted_sum[17] = $signed(-{in[0],2'b0})+$signed({in[25],1'b0})+$signed({in[1],1'b0})+$signed({in[10],1'b0})+$signed(-in[26])+$signed(in[28])+$signed(-{in[29],1'b0})+$signed(-in[5])+$signed(in[15])+$signed(sharing23_r)+$signed(-sharing24_r)+$signed(sharing34_r)+$signed(-1);
assign weighted_sum[18] = $signed(-{in[16],2'b0})+$signed(in[0])+$signed(-in[19])+$signed({in[4],1'b0})+$signed({in[30],1'b0})+$signed({in[31],2'b0})+$signed(sharing8_r)+$signed(-sharing9_r)+$signed(sharing35_r)+$signed(2);
assign weighted_sum[19] = $signed(-in[2])+$signed(-in[10])+$signed(-in[4])+$signed(-{in[13],1'b0})+$signed(-{in[22],1'b0})+$signed(sharing12_r)+$signed(sharing41_r)+$signed(-2);
assign weighted_sum[20] = $signed({in[16],2'b0})+$signed({in[8],1'b0})+$signed(in[24])+$signed(-{in[24],2'b0})+$signed(-{in[17],2'b0})+$signed(in[17])+$signed(-in[2])+$signed({in[3],2'b0})+$signed(in[27])+$signed({in[29],1'b0})+$signed({in[22],1'b0})+$signed(-{in[7],1'b0})+$signed(sharing13_r)+$signed(-sharing14_r)+$signed(sharing47_r)+$signed(-2);
assign weighted_sum[21] = $signed({in[22],2'b0})+$signed(-{in[8],1'b0})+$signed({in[10],1'b0})+$signed(-{in[18],1'b0})+$signed({in[27],1'b0})+$signed(in[11])+$signed({in[4],1'b0})+$signed({in[29],2'b0})+$signed(-{in[30],2'b0})+$signed(in[6])+$signed({in[23],1'b0})+$signed(sharing0_r)+$signed(-sharing1_r)+$signed(sharing38_r)+$signed(sharing47_r)+$signed(-1);
assign weighted_sum[22] = $signed(-{in[1],1'b0})+$signed({in[9],1'b0})+$signed(in[9])+$signed({in[26],2'b0})+$signed(in[10])+$signed({in[19],2'b0})+$signed({in[3],1'b0})+$signed(-{in[12],2'b0})+$signed(in[12])+$signed(-{in[13],2'b0})+$signed(in[29])+$signed({in[14],1'b0})+$signed(-in[31])+$signed(sharing19_r)+$signed(sharing20_r)+$signed(-sharing48_r)+$signed(2);
assign weighted_sum[23] = $signed(-{in[8],1'b0})+$signed(-in[0])+$signed(in[10])+$signed({in[12],1'b0})+$signed(-{in[29],1'b0})+$signed(-in[5])+$signed(-{in[30],3'b0})+$signed(in[6])+$signed(in[7])+$signed(sharing10_r)+$signed(-sharing11_r)+$signed(-sharing34_r)+$signed(sharing45_r)+$signed(0);
assign weighted_sum[24] = $signed(in[16])+$signed(-{in[17],2'b0})+$signed({in[25],1'b0})+$signed(-{in[10],1'b0})+$signed({in[3],1'b0})+$signed({in[29],1'b0})+$signed(-{in[6],2'b0})+$signed(in[30])+$signed(-{in[14],2'b0})+$signed(-in[23])+$signed(sharing21_r)+$signed(sharing22_r)+$signed(sharing36_r)+$signed(sharing37_r)+$signed(0);
assign weighted_sum[25] = $signed({in[8],1'b0})+$signed(in[25])+$signed(-{in[26],1'b0})+$signed(in[10])+$signed(-in[18])+$signed({in[20],1'b0})+$signed(-{in[29],2'b0})+$signed(-{in[13],1'b0})+$signed(in[30])+$signed({in[15],2'b0})+$signed(sharing23_r)+$signed(sharing24_r)+$signed(sharing38_r)+$signed(sharing48_r)+$signed(0);
assign weighted_sum[26] = $signed(-{in[24],2'b0})+$signed({in[16],1'b0})+$signed(in[25])+$signed(-in[17])+$signed(in[9])+$signed({in[3],2'b0})+$signed(-in[19])+$signed(in[4])+$signed(in[28])+$signed(-{in[5],1'b0})+$signed(in[13])+$signed(-in[21])+$signed(sharing25_r)+$signed(sharing26_r)+$signed(1);
assign weighted_sum[27] = $signed(in[22])+$signed(in[2])+$signed(-{in[19],1'b0})+$signed({in[3],1'b0})+$signed(-in[11])+$signed(-{in[20],2'b0})+$signed(in[4])+$signed({in[29],1'b0})+$signed({in[14],1'b0})+$signed(-in[30])+$signed(in[7])+$signed(-{in[15],2'b0})+$signed({in[7],1'b0})+$signed(in[23])+$signed(sharing27_r)+$signed(sharing28_r)+$signed(sharing39_r)+$signed(2);
assign weighted_sum[28] = $signed({in[8],1'b0})+$signed(-{in[25],2'b0})+$signed(-{in[27],2'b0})+$signed({in[19],1'b0})+$signed({in[12],1'b0})+$signed(-in[13])+$signed(-{in[15],1'b0})+$signed({in[23],1'b0})+$signed({in[30],1'b0})+$signed(-{in[31],1'b0})+$signed(sharing2_r)+$signed(-sharing3_r)+$signed(sharing40_r)+$signed(2);
assign weighted_sum[29] = $signed(in[16])+$signed(in[25])+$signed(-in[1])+$signed(-{in[2],2'b0})+$signed({in[18],1'b0})+$signed(in[2])+$signed({in[27],2'b0})+$signed({in[29],2'b0})+$signed(-{in[22],3'b0})+$signed(in[22])+$signed(sharing29_r)+$signed(sharing30_r)+$signed(-sharing39_r)+$signed(3);
assign weighted_sum[30] = $signed({in[8],2'b0})+$signed(-{in[16],1'b0})+$signed({in[22],1'b0})+$signed(-{in[17],1'b0})+$signed(-in[26])+$signed({in[11],1'b0})+$signed(in[29])+$signed(-{in[14],2'b0})+$signed({in[30],1'b0})+$signed({in[31],1'b0})+$signed(sharing27_r)+$signed(-sharing28_r)+$signed(-sharing43_r)+$signed(0);
assign weighted_sum[31] = $signed(-{in[16],2'b0})+$signed(in[16])+$signed({in[1],1'b0})+$signed(in[25])+$signed({in[18],1'b0})+$signed({in[26],1'b0})+$signed(-{in[19],2'b0})+$signed({in[11],1'b0})+$signed({in[28],2'b0})+$signed(in[4])+$signed(-{in[15],3'b0})+$signed({in[15],1'b0})+$signed(in[23])+$signed(sharing15_r)+$signed(-sharing16_r)+$signed(1);
assign out[0] = (weighted_sum[0][8]==1) ? 4'd0 : (weighted_sum[0][7:3] > 6 ? 4'd6 : weighted_sum[0][6:3]);
assign out[1] = (weighted_sum[1][8]==1) ? 4'd0 : (weighted_sum[1][7:3] > 6 ? 4'd6 : weighted_sum[1][6:3]);
assign out[2] = (weighted_sum[2][8]==1) ? 4'd0 : (weighted_sum[2][7:3] > 6 ? 4'd6 : weighted_sum[2][6:3]);
assign out[3] = (weighted_sum[3][8]==1) ? 4'd0 : (weighted_sum[3][7:3] > 6 ? 4'd6 : weighted_sum[3][6:3]);
assign out[4] = (weighted_sum[4][8]==1) ? 4'd0 : (weighted_sum[4][7:3] > 6 ? 4'd6 : weighted_sum[4][6:3]);
assign out[5] = (weighted_sum[5][8]==1) ? 4'd0 : (weighted_sum[5][7:3] > 6 ? 4'd6 : weighted_sum[5][6:3]);
assign out[6] = (weighted_sum[6][8]==1) ? 4'd0 : (weighted_sum[6][7:3] > 6 ? 4'd6 : weighted_sum[6][6:3]);
assign out[7] = (weighted_sum[7][8]==1) ? 4'd0 : (weighted_sum[7][7:3] > 6 ? 4'd6 : weighted_sum[7][6:3]);
assign out[8] = (weighted_sum[8][8]==1) ? 4'd0 : (weighted_sum[8][7:3] > 6 ? 4'd6 : weighted_sum[8][6:3]);
assign out[9] = (weighted_sum[9][8]==1) ? 4'd0 : (weighted_sum[9][7:3] > 6 ? 4'd6 : weighted_sum[9][6:3]);
assign out[10] = (weighted_sum[10][8]==1) ? 4'd0 : (weighted_sum[10][7:3] > 6 ? 4'd6 : weighted_sum[10][6:3]);
assign out[11] = (weighted_sum[11][8]==1) ? 4'd0 : (weighted_sum[11][7:3] > 6 ? 4'd6 : weighted_sum[11][6:3]);
assign out[12] = (weighted_sum[12][8]==1) ? 4'd0 : (weighted_sum[12][7:3] > 6 ? 4'd6 : weighted_sum[12][6:3]);
assign out[13] = (weighted_sum[13][8]==1) ? 4'd0 : (weighted_sum[13][7:3] > 6 ? 4'd6 : weighted_sum[13][6:3]);
assign out[14] = (weighted_sum[14][8]==1) ? 4'd0 : (weighted_sum[14][7:3] > 6 ? 4'd6 : weighted_sum[14][6:3]);
assign out[15] = (weighted_sum[15][8]==1) ? 4'd0 : (weighted_sum[15][7:3] > 6 ? 4'd6 : weighted_sum[15][6:3]);
assign out[16] = (weighted_sum[16][8]==1) ? 4'd0 : (weighted_sum[16][7:3] > 6 ? 4'd6 : weighted_sum[16][6:3]);
assign out[17] = (weighted_sum[17][8]==1) ? 4'd0 : (weighted_sum[17][7:3] > 6 ? 4'd6 : weighted_sum[17][6:3]);
assign out[18] = (weighted_sum[18][8]==1) ? 4'd0 : (weighted_sum[18][7:3] > 6 ? 4'd6 : weighted_sum[18][6:3]);
assign out[19] = (weighted_sum[19][8]==1) ? 4'd0 : (weighted_sum[19][7:3] > 6 ? 4'd6 : weighted_sum[19][6:3]);
assign out[20] = (weighted_sum[20][8]==1) ? 4'd0 : (weighted_sum[20][7:3] > 6 ? 4'd6 : weighted_sum[20][6:3]);
assign out[21] = (weighted_sum[21][8]==1) ? 4'd0 : (weighted_sum[21][7:3] > 6 ? 4'd6 : weighted_sum[21][6:3]);
assign out[22] = (weighted_sum[22][8]==1) ? 4'd0 : (weighted_sum[22][7:3] > 6 ? 4'd6 : weighted_sum[22][6:3]);
assign out[23] = (weighted_sum[23][8]==1) ? 4'd0 : (weighted_sum[23][7:3] > 6 ? 4'd6 : weighted_sum[23][6:3]);
assign out[24] = (weighted_sum[24][8]==1) ? 4'd0 : (weighted_sum[24][7:3] > 6 ? 4'd6 : weighted_sum[24][6:3]);
assign out[25] = (weighted_sum[25][8]==1) ? 4'd0 : (weighted_sum[25][7:3] > 6 ? 4'd6 : weighted_sum[25][6:3]);
assign out[26] = (weighted_sum[26][8]==1) ? 4'd0 : (weighted_sum[26][7:3] > 6 ? 4'd6 : weighted_sum[26][6:3]);
assign out[27] = (weighted_sum[27][8]==1) ? 4'd0 : (weighted_sum[27][7:3] > 6 ? 4'd6 : weighted_sum[27][6:3]);
assign out[28] = (weighted_sum[28][8]==1) ? 4'd0 : (weighted_sum[28][7:3] > 6 ? 4'd6 : weighted_sum[28][6:3]);
assign out[29] = (weighted_sum[29][8]==1) ? 4'd0 : (weighted_sum[29][7:3] > 6 ? 4'd6 : weighted_sum[29][6:3]);
assign out[30] = (weighted_sum[30][8]==1) ? 4'd0 : (weighted_sum[30][7:3] > 6 ? 4'd6 : weighted_sum[30][6:3]);
assign out[31] = (weighted_sum[31][8]==1) ? 4'd0 : (weighted_sum[31][7:3] > 6 ? 4'd6 : weighted_sum[31][6:3]);

always_ff @ (posedge clk or posedge rst) begin
	if (rst) begin
		sharing0_r <= 0;
		sharing1_r <= 0;
		sharing2_r <= 0;
		sharing3_r <= 0;
		sharing4_r <= 0;
		sharing5_r <= 0;
		sharing6_r <= 0;
		sharing7_r <= 0;
		sharing8_r <= 0;
		sharing9_r <= 0;
		sharing10_r <= 0;
		sharing11_r <= 0;
		sharing12_r <= 0;
		sharing13_r <= 0;
		sharing14_r <= 0;
		sharing15_r <= 0;
		sharing16_r <= 0;
		sharing17_r <= 0;
		sharing18_r <= 0;
		sharing19_r <= 0;
		sharing20_r <= 0;
		sharing21_r <= 0;
		sharing22_r <= 0;
		sharing23_r <= 0;
		sharing24_r <= 0;
		sharing25_r <= 0;
		sharing26_r <= 0;
		sharing27_r <= 0;
		sharing28_r <= 0;
		sharing29_r <= 0;
		sharing30_r <= 0;
		sharing31_r <= 0;
		sharing32_r <= 0;
		sharing33_r <= 0;
		sharing34_r <= 0;
		sharing35_r <= 0;
		sharing36_r <= 0;
		sharing37_r <= 0;
		sharing38_r <= 0;
		sharing39_r <= 0;
		sharing40_r <= 0;
		sharing41_r <= 0;
		sharing42_r <= 0;
		sharing43_r <= 0;
		sharing44_r <= 0;
		sharing45_r <= 0;
		sharing46_r <= 0;
		sharing47_r <= 0;
		sharing48_r <= 0;
		sharing49_r <= 0;
	end
	else begin
		sharing0_r <= sharing0_w;
		sharing1_r <= sharing1_w;
		sharing2_r <= sharing2_w;
		sharing3_r <= sharing3_w;
		sharing4_r <= sharing4_w;
		sharing5_r <= sharing5_w;
		sharing6_r <= sharing6_w;
		sharing7_r <= sharing7_w;
		sharing8_r <= sharing8_w;
		sharing9_r <= sharing9_w;
		sharing10_r <= sharing10_w;
		sharing11_r <= sharing11_w;
		sharing12_r <= sharing12_w;
		sharing13_r <= sharing13_w;
		sharing14_r <= sharing14_w;
		sharing15_r <= sharing15_w;
		sharing16_r <= sharing16_w;
		sharing17_r <= sharing17_w;
		sharing18_r <= sharing18_w;
		sharing19_r <= sharing19_w;
		sharing20_r <= sharing20_w;
		sharing21_r <= sharing21_w;
		sharing22_r <= sharing22_w;
		sharing23_r <= sharing23_w;
		sharing24_r <= sharing24_w;
		sharing25_r <= sharing25_w;
		sharing26_r <= sharing26_w;
		sharing27_r <= sharing27_w;
		sharing28_r <= sharing28_w;
		sharing29_r <= sharing29_w;
		sharing30_r <= sharing30_w;
		sharing31_r <= sharing31_w;
		sharing32_r <= sharing32_w;
		sharing33_r <= sharing33_w;
		sharing34_r <= sharing34_w;
		sharing35_r <= sharing35_w;
		sharing36_r <= sharing36_w;
		sharing37_r <= sharing37_w;
		sharing38_r <= sharing38_w;
		sharing39_r <= sharing39_w;
		sharing40_r <= sharing40_w;
		sharing41_r <= sharing41_w;
		sharing42_r <= sharing42_w;
		sharing43_r <= sharing43_w;
		sharing44_r <= sharing44_w;
		sharing45_r <= sharing45_w;
		sharing46_r <= sharing46_w;
		sharing47_r <= sharing47_w;
		sharing48_r <= sharing48_w;
		sharing49_r <= sharing49_w;
	end
end
endmodule
